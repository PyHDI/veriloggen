

module top
(
  input clk,
  input btnCpuReset,
  input btnC,
  input btnU,
  input btnL,
  input btnR,
  input btnD,
  input [16-1:0] sw,
  output [16-1:0] led
);

  wire new_CLK;
  assign new_CLK = clk;
  reg RST_X;
  reg RST;

  always @(posedge clk) begin
    RST_X <= btnCpuReset;
    RST <= !RST_X;
  end


  blinkled
  inst_blinkled
  (
    .CLK(new_CLK),
    .RST(RST),
    .btnC(btnC),
    .btnU(btnU),
    .btnL(btnL),
    .btnR(btnR),
    .btnD(btnD),
    .sw(sw),
    .led(led)
  );


endmodule



module blinkled
(
  input CLK,
  input RST,
  input btnC,
  input btnU,
  input btnL,
  input btnR,
  input btnD,
  input [16-1:0] sw,
  output [16-1:0] led
);

  reg [15-1:0] count;
  reg done;
  assign led = { done, count };
  reg _mymutex_lock_reg;
  reg [32-1:0] _mymutex_lock_id;
  reg [64-1:0] _th_myfunc_start;
  reg [32-1:0] th_blink;
  localparam th_blink_init = 0;
  reg signed [32-1:0] _th_blink_polarity_259;
  reg signed [32-1:0] _th_blink_tid_260;
  reg [32-1:0] th_myfunc_0;
  localparam th_myfunc_0_init = 0;
  reg [32-1:0] th_myfunc_1;
  localparam th_myfunc_1_init = 0;
  reg [32-1:0] th_myfunc_2;
  localparam th_myfunc_2_init = 0;
  reg [32-1:0] th_myfunc_3;
  localparam th_myfunc_3_init = 0;
  reg [32-1:0] th_myfunc_4;
  localparam th_myfunc_4_init = 0;
  reg [32-1:0] th_myfunc_5;
  localparam th_myfunc_5_init = 0;
  reg [32-1:0] th_myfunc_6;
  localparam th_myfunc_6_init = 0;
  reg [32-1:0] th_myfunc_7;
  localparam th_myfunc_7_init = 0;
  reg [32-1:0] th_myfunc_8;
  localparam th_myfunc_8_init = 0;
  reg [32-1:0] th_myfunc_9;
  localparam th_myfunc_9_init = 0;
  reg [32-1:0] th_myfunc_10;
  localparam th_myfunc_10_init = 0;
  reg [32-1:0] th_myfunc_11;
  localparam th_myfunc_11_init = 0;
  reg [32-1:0] th_myfunc_12;
  localparam th_myfunc_12_init = 0;
  reg [32-1:0] th_myfunc_13;
  localparam th_myfunc_13_init = 0;
  reg [32-1:0] th_myfunc_14;
  localparam th_myfunc_14_init = 0;
  reg [32-1:0] th_myfunc_15;
  localparam th_myfunc_15_init = 0;
  reg [32-1:0] th_myfunc_16;
  localparam th_myfunc_16_init = 0;
  reg [32-1:0] th_myfunc_17;
  localparam th_myfunc_17_init = 0;
  reg [32-1:0] th_myfunc_18;
  localparam th_myfunc_18_init = 0;
  reg [32-1:0] th_myfunc_19;
  localparam th_myfunc_19_init = 0;
  reg [32-1:0] th_myfunc_20;
  localparam th_myfunc_20_init = 0;
  reg [32-1:0] th_myfunc_21;
  localparam th_myfunc_21_init = 0;
  reg [32-1:0] th_myfunc_22;
  localparam th_myfunc_22_init = 0;
  reg [32-1:0] th_myfunc_23;
  localparam th_myfunc_23_init = 0;
  reg [32-1:0] th_myfunc_24;
  localparam th_myfunc_24_init = 0;
  reg [32-1:0] th_myfunc_25;
  localparam th_myfunc_25_init = 0;
  reg [32-1:0] th_myfunc_26;
  localparam th_myfunc_26_init = 0;
  reg [32-1:0] th_myfunc_27;
  localparam th_myfunc_27_init = 0;
  reg [32-1:0] th_myfunc_28;
  localparam th_myfunc_28_init = 0;
  reg [32-1:0] th_myfunc_29;
  localparam th_myfunc_29_init = 0;
  reg [32-1:0] th_myfunc_30;
  localparam th_myfunc_30_init = 0;
  reg [32-1:0] th_myfunc_31;
  localparam th_myfunc_31_init = 0;
  reg [32-1:0] th_myfunc_32;
  localparam th_myfunc_32_init = 0;
  reg [32-1:0] th_myfunc_33;
  localparam th_myfunc_33_init = 0;
  reg [32-1:0] th_myfunc_34;
  localparam th_myfunc_34_init = 0;
  reg [32-1:0] th_myfunc_35;
  localparam th_myfunc_35_init = 0;
  reg [32-1:0] th_myfunc_36;
  localparam th_myfunc_36_init = 0;
  reg [32-1:0] th_myfunc_37;
  localparam th_myfunc_37_init = 0;
  reg [32-1:0] th_myfunc_38;
  localparam th_myfunc_38_init = 0;
  reg [32-1:0] th_myfunc_39;
  localparam th_myfunc_39_init = 0;
  reg [32-1:0] th_myfunc_40;
  localparam th_myfunc_40_init = 0;
  reg [32-1:0] th_myfunc_41;
  localparam th_myfunc_41_init = 0;
  reg [32-1:0] th_myfunc_42;
  localparam th_myfunc_42_init = 0;
  reg [32-1:0] th_myfunc_43;
  localparam th_myfunc_43_init = 0;
  reg [32-1:0] th_myfunc_44;
  localparam th_myfunc_44_init = 0;
  reg [32-1:0] th_myfunc_45;
  localparam th_myfunc_45_init = 0;
  reg [32-1:0] th_myfunc_46;
  localparam th_myfunc_46_init = 0;
  reg [32-1:0] th_myfunc_47;
  localparam th_myfunc_47_init = 0;
  reg [32-1:0] th_myfunc_48;
  localparam th_myfunc_48_init = 0;
  reg [32-1:0] th_myfunc_49;
  localparam th_myfunc_49_init = 0;
  reg [32-1:0] th_myfunc_50;
  localparam th_myfunc_50_init = 0;
  reg [32-1:0] th_myfunc_51;
  localparam th_myfunc_51_init = 0;
  reg [32-1:0] th_myfunc_52;
  localparam th_myfunc_52_init = 0;
  reg [32-1:0] th_myfunc_53;
  localparam th_myfunc_53_init = 0;
  reg [32-1:0] th_myfunc_54;
  localparam th_myfunc_54_init = 0;
  reg [32-1:0] th_myfunc_55;
  localparam th_myfunc_55_init = 0;
  reg [32-1:0] th_myfunc_56;
  localparam th_myfunc_56_init = 0;
  reg [32-1:0] th_myfunc_57;
  localparam th_myfunc_57_init = 0;
  reg [32-1:0] th_myfunc_58;
  localparam th_myfunc_58_init = 0;
  reg [32-1:0] th_myfunc_59;
  localparam th_myfunc_59_init = 0;
  reg [32-1:0] th_myfunc_60;
  localparam th_myfunc_60_init = 0;
  reg [32-1:0] th_myfunc_61;
  localparam th_myfunc_61_init = 0;
  reg [32-1:0] th_myfunc_62;
  localparam th_myfunc_62_init = 0;
  reg [32-1:0] th_myfunc_63;
  localparam th_myfunc_63_init = 0;
  reg _th_myfunc_0_called;
  reg signed [32-1:0] _th_myfunc_0_tid_261;
  reg signed [32-1:0] _th_myfunc_0_tid_262;
  reg signed [32-1:0] _th_myfunc_0_time_263;
  reg signed [32-1:0] _th_myfunc_0_i_264;
  reg _th_myfunc_1_called;
  reg signed [32-1:0] _th_myfunc_1_tid_265;
  reg signed [32-1:0] _th_myfunc_1_tid_266;
  reg signed [32-1:0] _th_myfunc_1_time_267;
  reg signed [32-1:0] _th_myfunc_1_i_268;
  reg _th_myfunc_2_called;
  reg signed [32-1:0] _th_myfunc_2_tid_269;
  reg signed [32-1:0] _th_myfunc_2_tid_270;
  reg signed [32-1:0] _th_myfunc_2_time_271;
  reg signed [32-1:0] _th_myfunc_2_i_272;
  reg _th_myfunc_3_called;
  reg signed [32-1:0] _th_myfunc_3_tid_273;
  reg signed [32-1:0] _th_myfunc_3_tid_274;
  reg signed [32-1:0] _th_myfunc_3_time_275;
  reg signed [32-1:0] _th_myfunc_3_i_276;
  reg _th_myfunc_4_called;
  reg signed [32-1:0] _th_myfunc_4_tid_277;
  reg signed [32-1:0] _th_myfunc_4_tid_278;
  reg signed [32-1:0] _th_myfunc_4_time_279;
  reg signed [32-1:0] _th_myfunc_4_i_280;
  reg _th_myfunc_5_called;
  reg signed [32-1:0] _th_myfunc_5_tid_281;
  reg signed [32-1:0] _th_myfunc_5_tid_282;
  reg signed [32-1:0] _th_myfunc_5_time_283;
  reg signed [32-1:0] _th_myfunc_5_i_284;
  reg _th_myfunc_6_called;
  reg signed [32-1:0] _th_myfunc_6_tid_285;
  reg signed [32-1:0] _th_myfunc_6_tid_286;
  reg signed [32-1:0] _th_myfunc_6_time_287;
  reg signed [32-1:0] _th_myfunc_6_i_288;
  reg _th_myfunc_7_called;
  reg signed [32-1:0] _th_myfunc_7_tid_289;
  reg signed [32-1:0] _th_myfunc_7_tid_290;
  reg signed [32-1:0] _th_myfunc_7_time_291;
  reg signed [32-1:0] _th_myfunc_7_i_292;
  reg _th_myfunc_8_called;
  reg signed [32-1:0] _th_myfunc_8_tid_293;
  reg signed [32-1:0] _th_myfunc_8_tid_294;
  reg signed [32-1:0] _th_myfunc_8_time_295;
  reg signed [32-1:0] _th_myfunc_8_i_296;
  reg _th_myfunc_9_called;
  reg signed [32-1:0] _th_myfunc_9_tid_297;
  reg signed [32-1:0] _th_myfunc_9_tid_298;
  reg signed [32-1:0] _th_myfunc_9_time_299;
  reg signed [32-1:0] _th_myfunc_9_i_300;
  reg _th_myfunc_10_called;
  reg signed [32-1:0] _th_myfunc_10_tid_301;
  reg signed [32-1:0] _th_myfunc_10_tid_302;
  reg signed [32-1:0] _th_myfunc_10_time_303;
  reg signed [32-1:0] _th_myfunc_10_i_304;
  reg _th_myfunc_11_called;
  reg signed [32-1:0] _th_myfunc_11_tid_305;
  reg signed [32-1:0] _th_myfunc_11_tid_306;
  reg signed [32-1:0] _th_myfunc_11_time_307;
  reg signed [32-1:0] _th_myfunc_11_i_308;
  reg _th_myfunc_12_called;
  reg signed [32-1:0] _th_myfunc_12_tid_309;
  reg signed [32-1:0] _th_myfunc_12_tid_310;
  reg signed [32-1:0] _th_myfunc_12_time_311;
  reg signed [32-1:0] _th_myfunc_12_i_312;
  reg _th_myfunc_13_called;
  reg signed [32-1:0] _th_myfunc_13_tid_313;
  reg signed [32-1:0] _th_myfunc_13_tid_314;
  reg signed [32-1:0] _th_myfunc_13_time_315;
  reg signed [32-1:0] _th_myfunc_13_i_316;
  reg _th_myfunc_14_called;
  reg signed [32-1:0] _th_myfunc_14_tid_317;
  reg signed [32-1:0] _th_myfunc_14_tid_318;
  reg signed [32-1:0] _th_myfunc_14_time_319;
  reg signed [32-1:0] _th_myfunc_14_i_320;
  reg _th_myfunc_15_called;
  reg signed [32-1:0] _th_myfunc_15_tid_321;
  reg signed [32-1:0] _th_myfunc_15_tid_322;
  reg signed [32-1:0] _th_myfunc_15_time_323;
  reg signed [32-1:0] _th_myfunc_15_i_324;
  reg _th_myfunc_16_called;
  reg signed [32-1:0] _th_myfunc_16_tid_325;
  reg signed [32-1:0] _th_myfunc_16_tid_326;
  reg signed [32-1:0] _th_myfunc_16_time_327;
  reg signed [32-1:0] _th_myfunc_16_i_328;
  reg _th_myfunc_17_called;
  reg signed [32-1:0] _th_myfunc_17_tid_329;
  reg signed [32-1:0] _th_myfunc_17_tid_330;
  reg signed [32-1:0] _th_myfunc_17_time_331;
  reg signed [32-1:0] _th_myfunc_17_i_332;
  reg _th_myfunc_18_called;
  reg signed [32-1:0] _th_myfunc_18_tid_333;
  reg signed [32-1:0] _th_myfunc_18_tid_334;
  reg signed [32-1:0] _th_myfunc_18_time_335;
  reg signed [32-1:0] _th_myfunc_18_i_336;
  reg _th_myfunc_19_called;
  reg signed [32-1:0] _th_myfunc_19_tid_337;
  reg signed [32-1:0] _th_myfunc_19_tid_338;
  reg signed [32-1:0] _th_myfunc_19_time_339;
  reg signed [32-1:0] _th_myfunc_19_i_340;
  reg _th_myfunc_20_called;
  reg signed [32-1:0] _th_myfunc_20_tid_341;
  reg signed [32-1:0] _th_myfunc_20_tid_342;
  reg signed [32-1:0] _th_myfunc_20_time_343;
  reg signed [32-1:0] _th_myfunc_20_i_344;
  reg _th_myfunc_21_called;
  reg signed [32-1:0] _th_myfunc_21_tid_345;
  reg signed [32-1:0] _th_myfunc_21_tid_346;
  reg signed [32-1:0] _th_myfunc_21_time_347;
  reg signed [32-1:0] _th_myfunc_21_i_348;
  reg _th_myfunc_22_called;
  reg signed [32-1:0] _th_myfunc_22_tid_349;
  reg signed [32-1:0] _th_myfunc_22_tid_350;
  reg signed [32-1:0] _th_myfunc_22_time_351;
  reg signed [32-1:0] _th_myfunc_22_i_352;
  reg _th_myfunc_23_called;
  reg signed [32-1:0] _th_myfunc_23_tid_353;
  reg signed [32-1:0] _th_myfunc_23_tid_354;
  reg signed [32-1:0] _th_myfunc_23_time_355;
  reg signed [32-1:0] _th_myfunc_23_i_356;
  reg _th_myfunc_24_called;
  reg signed [32-1:0] _th_myfunc_24_tid_357;
  reg signed [32-1:0] _th_myfunc_24_tid_358;
  reg signed [32-1:0] _th_myfunc_24_time_359;
  reg signed [32-1:0] _th_myfunc_24_i_360;
  reg _th_myfunc_25_called;
  reg signed [32-1:0] _th_myfunc_25_tid_361;
  reg signed [32-1:0] _th_myfunc_25_tid_362;
  reg signed [32-1:0] _th_myfunc_25_time_363;
  reg signed [32-1:0] _th_myfunc_25_i_364;
  reg _th_myfunc_26_called;
  reg signed [32-1:0] _th_myfunc_26_tid_365;
  reg signed [32-1:0] _th_myfunc_26_tid_366;
  reg signed [32-1:0] _th_myfunc_26_time_367;
  reg signed [32-1:0] _th_myfunc_26_i_368;
  reg _th_myfunc_27_called;
  reg signed [32-1:0] _th_myfunc_27_tid_369;
  reg signed [32-1:0] _th_myfunc_27_tid_370;
  reg signed [32-1:0] _th_myfunc_27_time_371;
  reg signed [32-1:0] _th_myfunc_27_i_372;
  reg _th_myfunc_28_called;
  reg signed [32-1:0] _th_myfunc_28_tid_373;
  reg signed [32-1:0] _th_myfunc_28_tid_374;
  reg signed [32-1:0] _th_myfunc_28_time_375;
  reg signed [32-1:0] _th_myfunc_28_i_376;
  reg _th_myfunc_29_called;
  reg signed [32-1:0] _th_myfunc_29_tid_377;
  reg signed [32-1:0] _th_myfunc_29_tid_378;
  reg signed [32-1:0] _th_myfunc_29_time_379;
  reg signed [32-1:0] _th_myfunc_29_i_380;
  reg _th_myfunc_30_called;
  reg signed [32-1:0] _th_myfunc_30_tid_381;
  reg signed [32-1:0] _th_myfunc_30_tid_382;
  reg signed [32-1:0] _th_myfunc_30_time_383;
  reg signed [32-1:0] _th_myfunc_30_i_384;
  reg _th_myfunc_31_called;
  reg signed [32-1:0] _th_myfunc_31_tid_385;
  reg signed [32-1:0] _th_myfunc_31_tid_386;
  reg signed [32-1:0] _th_myfunc_31_time_387;
  reg signed [32-1:0] _th_myfunc_31_i_388;
  reg _th_myfunc_32_called;
  reg signed [32-1:0] _th_myfunc_32_tid_389;
  reg signed [32-1:0] _th_myfunc_32_tid_390;
  reg signed [32-1:0] _th_myfunc_32_time_391;
  reg signed [32-1:0] _th_myfunc_32_i_392;
  reg _th_myfunc_33_called;
  reg signed [32-1:0] _th_myfunc_33_tid_393;
  reg signed [32-1:0] _th_myfunc_33_tid_394;
  reg signed [32-1:0] _th_myfunc_33_time_395;
  reg signed [32-1:0] _th_myfunc_33_i_396;
  reg _th_myfunc_34_called;
  reg signed [32-1:0] _th_myfunc_34_tid_397;
  reg signed [32-1:0] _th_myfunc_34_tid_398;
  reg signed [32-1:0] _th_myfunc_34_time_399;
  reg signed [32-1:0] _th_myfunc_34_i_400;
  reg _th_myfunc_35_called;
  reg signed [32-1:0] _th_myfunc_35_tid_401;
  reg signed [32-1:0] _th_myfunc_35_tid_402;
  reg signed [32-1:0] _th_myfunc_35_time_403;
  reg signed [32-1:0] _th_myfunc_35_i_404;
  reg _th_myfunc_36_called;
  reg signed [32-1:0] _th_myfunc_36_tid_405;
  reg signed [32-1:0] _th_myfunc_36_tid_406;
  reg signed [32-1:0] _th_myfunc_36_time_407;
  reg signed [32-1:0] _th_myfunc_36_i_408;
  reg _th_myfunc_37_called;
  reg signed [32-1:0] _th_myfunc_37_tid_409;
  reg signed [32-1:0] _th_myfunc_37_tid_410;
  reg signed [32-1:0] _th_myfunc_37_time_411;
  reg signed [32-1:0] _th_myfunc_37_i_412;
  reg _th_myfunc_38_called;
  reg signed [32-1:0] _th_myfunc_38_tid_413;
  reg signed [32-1:0] _th_myfunc_38_tid_414;
  reg signed [32-1:0] _th_myfunc_38_time_415;
  reg signed [32-1:0] _th_myfunc_38_i_416;
  reg _th_myfunc_39_called;
  reg signed [32-1:0] _th_myfunc_39_tid_417;
  reg signed [32-1:0] _th_myfunc_39_tid_418;
  reg signed [32-1:0] _th_myfunc_39_time_419;
  reg signed [32-1:0] _th_myfunc_39_i_420;
  reg _th_myfunc_40_called;
  reg signed [32-1:0] _th_myfunc_40_tid_421;
  reg signed [32-1:0] _th_myfunc_40_tid_422;
  reg signed [32-1:0] _th_myfunc_40_time_423;
  reg signed [32-1:0] _th_myfunc_40_i_424;
  reg _th_myfunc_41_called;
  reg signed [32-1:0] _th_myfunc_41_tid_425;
  reg signed [32-1:0] _th_myfunc_41_tid_426;
  reg signed [32-1:0] _th_myfunc_41_time_427;
  reg signed [32-1:0] _th_myfunc_41_i_428;
  reg _th_myfunc_42_called;
  reg signed [32-1:0] _th_myfunc_42_tid_429;
  reg signed [32-1:0] _th_myfunc_42_tid_430;
  reg signed [32-1:0] _th_myfunc_42_time_431;
  reg signed [32-1:0] _th_myfunc_42_i_432;
  reg _th_myfunc_43_called;
  reg signed [32-1:0] _th_myfunc_43_tid_433;
  reg signed [32-1:0] _th_myfunc_43_tid_434;
  reg signed [32-1:0] _th_myfunc_43_time_435;
  reg signed [32-1:0] _th_myfunc_43_i_436;
  reg _th_myfunc_44_called;
  reg signed [32-1:0] _th_myfunc_44_tid_437;
  reg signed [32-1:0] _th_myfunc_44_tid_438;
  reg signed [32-1:0] _th_myfunc_44_time_439;
  reg signed [32-1:0] _th_myfunc_44_i_440;
  reg _th_myfunc_45_called;
  reg signed [32-1:0] _th_myfunc_45_tid_441;
  reg signed [32-1:0] _th_myfunc_45_tid_442;
  reg signed [32-1:0] _th_myfunc_45_time_443;
  reg signed [32-1:0] _th_myfunc_45_i_444;
  reg _th_myfunc_46_called;
  reg signed [32-1:0] _th_myfunc_46_tid_445;
  reg signed [32-1:0] _th_myfunc_46_tid_446;
  reg signed [32-1:0] _th_myfunc_46_time_447;
  reg signed [32-1:0] _th_myfunc_46_i_448;
  reg _th_myfunc_47_called;
  reg signed [32-1:0] _th_myfunc_47_tid_449;
  reg signed [32-1:0] _th_myfunc_47_tid_450;
  reg signed [32-1:0] _th_myfunc_47_time_451;
  reg signed [32-1:0] _th_myfunc_47_i_452;
  reg _th_myfunc_48_called;
  reg signed [32-1:0] _th_myfunc_48_tid_453;
  reg signed [32-1:0] _th_myfunc_48_tid_454;
  reg signed [32-1:0] _th_myfunc_48_time_455;
  reg signed [32-1:0] _th_myfunc_48_i_456;
  reg _th_myfunc_49_called;
  reg signed [32-1:0] _th_myfunc_49_tid_457;
  reg signed [32-1:0] _th_myfunc_49_tid_458;
  reg signed [32-1:0] _th_myfunc_49_time_459;
  reg signed [32-1:0] _th_myfunc_49_i_460;
  reg _th_myfunc_50_called;
  reg signed [32-1:0] _th_myfunc_50_tid_461;
  reg signed [32-1:0] _th_myfunc_50_tid_462;
  reg signed [32-1:0] _th_myfunc_50_time_463;
  reg signed [32-1:0] _th_myfunc_50_i_464;
  reg _th_myfunc_51_called;
  reg signed [32-1:0] _th_myfunc_51_tid_465;
  reg signed [32-1:0] _th_myfunc_51_tid_466;
  reg signed [32-1:0] _th_myfunc_51_time_467;
  reg signed [32-1:0] _th_myfunc_51_i_468;
  reg _th_myfunc_52_called;
  reg signed [32-1:0] _th_myfunc_52_tid_469;
  reg signed [32-1:0] _th_myfunc_52_tid_470;
  reg signed [32-1:0] _th_myfunc_52_time_471;
  reg signed [32-1:0] _th_myfunc_52_i_472;
  reg _th_myfunc_53_called;
  reg signed [32-1:0] _th_myfunc_53_tid_473;
  reg signed [32-1:0] _th_myfunc_53_tid_474;
  reg signed [32-1:0] _th_myfunc_53_time_475;
  reg signed [32-1:0] _th_myfunc_53_i_476;
  reg _th_myfunc_54_called;
  reg signed [32-1:0] _th_myfunc_54_tid_477;
  reg signed [32-1:0] _th_myfunc_54_tid_478;
  reg signed [32-1:0] _th_myfunc_54_time_479;
  reg signed [32-1:0] _th_myfunc_54_i_480;
  reg _th_myfunc_55_called;
  reg signed [32-1:0] _th_myfunc_55_tid_481;
  reg signed [32-1:0] _th_myfunc_55_tid_482;
  reg signed [32-1:0] _th_myfunc_55_time_483;
  reg signed [32-1:0] _th_myfunc_55_i_484;
  reg _th_myfunc_56_called;
  reg signed [32-1:0] _th_myfunc_56_tid_485;
  reg signed [32-1:0] _th_myfunc_56_tid_486;
  reg signed [32-1:0] _th_myfunc_56_time_487;
  reg signed [32-1:0] _th_myfunc_56_i_488;
  reg _th_myfunc_57_called;
  reg signed [32-1:0] _th_myfunc_57_tid_489;
  reg signed [32-1:0] _th_myfunc_57_tid_490;
  reg signed [32-1:0] _th_myfunc_57_time_491;
  reg signed [32-1:0] _th_myfunc_57_i_492;
  reg _th_myfunc_58_called;
  reg signed [32-1:0] _th_myfunc_58_tid_493;
  reg signed [32-1:0] _th_myfunc_58_tid_494;
  reg signed [32-1:0] _th_myfunc_58_time_495;
  reg signed [32-1:0] _th_myfunc_58_i_496;
  reg _th_myfunc_59_called;
  reg signed [32-1:0] _th_myfunc_59_tid_497;
  reg signed [32-1:0] _th_myfunc_59_tid_498;
  reg signed [32-1:0] _th_myfunc_59_time_499;
  reg signed [32-1:0] _th_myfunc_59_i_500;
  reg _th_myfunc_60_called;
  reg signed [32-1:0] _th_myfunc_60_tid_501;
  reg signed [32-1:0] _th_myfunc_60_tid_502;
  reg signed [32-1:0] _th_myfunc_60_time_503;
  reg signed [32-1:0] _th_myfunc_60_i_504;
  reg _th_myfunc_61_called;
  reg signed [32-1:0] _th_myfunc_61_tid_505;
  reg signed [32-1:0] _th_myfunc_61_tid_506;
  reg signed [32-1:0] _th_myfunc_61_time_507;
  reg signed [32-1:0] _th_myfunc_61_i_508;
  reg _th_myfunc_62_called;
  reg signed [32-1:0] _th_myfunc_62_tid_509;
  reg signed [32-1:0] _th_myfunc_62_tid_510;
  reg signed [32-1:0] _th_myfunc_62_time_511;
  reg signed [32-1:0] _th_myfunc_62_i_512;
  reg _th_myfunc_63_called;
  reg signed [32-1:0] _th_myfunc_63_tid_513;
  reg signed [32-1:0] _th_myfunc_63_tid_514;
  reg signed [32-1:0] _th_myfunc_63_time_515;
  reg signed [32-1:0] _th_myfunc_63_i_516;

  always @(posedge CLK) begin
    if(RST) begin
      _mymutex_lock_reg <= 0;
      _mymutex_lock_id <= 0;
    end else begin
      if((th_myfunc_0 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 0;
      end 
      if((th_myfunc_0 == 11) && (_mymutex_lock_id == 0)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_1 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 1;
      end 
      if((th_myfunc_1 == 11) && (_mymutex_lock_id == 1)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_2 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 2;
      end 
      if((th_myfunc_2 == 11) && (_mymutex_lock_id == 2)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_3 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 3;
      end 
      if((th_myfunc_3 == 11) && (_mymutex_lock_id == 3)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_4 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 4;
      end 
      if((th_myfunc_4 == 11) && (_mymutex_lock_id == 4)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_5 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 5;
      end 
      if((th_myfunc_5 == 11) && (_mymutex_lock_id == 5)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_6 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 6;
      end 
      if((th_myfunc_6 == 11) && (_mymutex_lock_id == 6)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_7 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 7;
      end 
      if((th_myfunc_7 == 11) && (_mymutex_lock_id == 7)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_8 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 8;
      end 
      if((th_myfunc_8 == 11) && (_mymutex_lock_id == 8)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_9 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 9;
      end 
      if((th_myfunc_9 == 11) && (_mymutex_lock_id == 9)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_10 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 10;
      end 
      if((th_myfunc_10 == 11) && (_mymutex_lock_id == 10)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_11 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 11;
      end 
      if((th_myfunc_11 == 11) && (_mymutex_lock_id == 11)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_12 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 12;
      end 
      if((th_myfunc_12 == 11) && (_mymutex_lock_id == 12)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_13 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 13;
      end 
      if((th_myfunc_13 == 11) && (_mymutex_lock_id == 13)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_14 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 14;
      end 
      if((th_myfunc_14 == 11) && (_mymutex_lock_id == 14)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_15 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 15;
      end 
      if((th_myfunc_15 == 11) && (_mymutex_lock_id == 15)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_16 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 16;
      end 
      if((th_myfunc_16 == 11) && (_mymutex_lock_id == 16)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_17 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 17;
      end 
      if((th_myfunc_17 == 11) && (_mymutex_lock_id == 17)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_18 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 18;
      end 
      if((th_myfunc_18 == 11) && (_mymutex_lock_id == 18)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_19 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 19;
      end 
      if((th_myfunc_19 == 11) && (_mymutex_lock_id == 19)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_20 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 20;
      end 
      if((th_myfunc_20 == 11) && (_mymutex_lock_id == 20)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_21 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 21;
      end 
      if((th_myfunc_21 == 11) && (_mymutex_lock_id == 21)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_22 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 22;
      end 
      if((th_myfunc_22 == 11) && (_mymutex_lock_id == 22)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_23 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 23;
      end 
      if((th_myfunc_23 == 11) && (_mymutex_lock_id == 23)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_24 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 24;
      end 
      if((th_myfunc_24 == 11) && (_mymutex_lock_id == 24)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_25 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 25;
      end 
      if((th_myfunc_25 == 11) && (_mymutex_lock_id == 25)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_26 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 26;
      end 
      if((th_myfunc_26 == 11) && (_mymutex_lock_id == 26)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_27 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 27;
      end 
      if((th_myfunc_27 == 11) && (_mymutex_lock_id == 27)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_28 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 28;
      end 
      if((th_myfunc_28 == 11) && (_mymutex_lock_id == 28)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_29 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 29;
      end 
      if((th_myfunc_29 == 11) && (_mymutex_lock_id == 29)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_30 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 30;
      end 
      if((th_myfunc_30 == 11) && (_mymutex_lock_id == 30)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_31 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 31;
      end 
      if((th_myfunc_31 == 11) && (_mymutex_lock_id == 31)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_32 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 32;
      end 
      if((th_myfunc_32 == 11) && (_mymutex_lock_id == 32)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_33 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 33;
      end 
      if((th_myfunc_33 == 11) && (_mymutex_lock_id == 33)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_34 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 34;
      end 
      if((th_myfunc_34 == 11) && (_mymutex_lock_id == 34)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_35 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 35;
      end 
      if((th_myfunc_35 == 11) && (_mymutex_lock_id == 35)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_36 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 36;
      end 
      if((th_myfunc_36 == 11) && (_mymutex_lock_id == 36)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_37 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 37;
      end 
      if((th_myfunc_37 == 11) && (_mymutex_lock_id == 37)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_38 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 38;
      end 
      if((th_myfunc_38 == 11) && (_mymutex_lock_id == 38)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_39 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 39;
      end 
      if((th_myfunc_39 == 11) && (_mymutex_lock_id == 39)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_40 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 40;
      end 
      if((th_myfunc_40 == 11) && (_mymutex_lock_id == 40)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_41 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 41;
      end 
      if((th_myfunc_41 == 11) && (_mymutex_lock_id == 41)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_42 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 42;
      end 
      if((th_myfunc_42 == 11) && (_mymutex_lock_id == 42)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_43 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 43;
      end 
      if((th_myfunc_43 == 11) && (_mymutex_lock_id == 43)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_44 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 44;
      end 
      if((th_myfunc_44 == 11) && (_mymutex_lock_id == 44)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_45 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 45;
      end 
      if((th_myfunc_45 == 11) && (_mymutex_lock_id == 45)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_46 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 46;
      end 
      if((th_myfunc_46 == 11) && (_mymutex_lock_id == 46)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_47 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 47;
      end 
      if((th_myfunc_47 == 11) && (_mymutex_lock_id == 47)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_48 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 48;
      end 
      if((th_myfunc_48 == 11) && (_mymutex_lock_id == 48)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_49 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 49;
      end 
      if((th_myfunc_49 == 11) && (_mymutex_lock_id == 49)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_50 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 50;
      end 
      if((th_myfunc_50 == 11) && (_mymutex_lock_id == 50)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_51 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 51;
      end 
      if((th_myfunc_51 == 11) && (_mymutex_lock_id == 51)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_52 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 52;
      end 
      if((th_myfunc_52 == 11) && (_mymutex_lock_id == 52)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_53 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 53;
      end 
      if((th_myfunc_53 == 11) && (_mymutex_lock_id == 53)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_54 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 54;
      end 
      if((th_myfunc_54 == 11) && (_mymutex_lock_id == 54)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_55 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 55;
      end 
      if((th_myfunc_55 == 11) && (_mymutex_lock_id == 55)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_56 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 56;
      end 
      if((th_myfunc_56 == 11) && (_mymutex_lock_id == 56)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_57 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 57;
      end 
      if((th_myfunc_57 == 11) && (_mymutex_lock_id == 57)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_58 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 58;
      end 
      if((th_myfunc_58 == 11) && (_mymutex_lock_id == 58)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_59 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 59;
      end 
      if((th_myfunc_59 == 11) && (_mymutex_lock_id == 59)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_60 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 60;
      end 
      if((th_myfunc_60 == 11) && (_mymutex_lock_id == 60)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_61 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 61;
      end 
      if((th_myfunc_61 == 11) && (_mymutex_lock_id == 61)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_62 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 62;
      end 
      if((th_myfunc_62 == 11) && (_mymutex_lock_id == 62)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_63 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 63;
      end 
      if((th_myfunc_63 == 11) && (_mymutex_lock_id == 63)) begin
        _mymutex_lock_reg <= 0;
      end 
    end
  end

  localparam th_blink_1 = 1;
  localparam th_blink_2 = 2;
  localparam th_blink_3 = 3;
  localparam th_blink_4 = 4;
  localparam th_blink_5 = 5;
  localparam th_blink_6 = 6;
  localparam th_blink_7 = 7;
  localparam th_blink_8 = 8;
  localparam th_blink_9 = 9;
  localparam th_blink_10 = 10;
  localparam th_blink_11 = 11;
  localparam th_blink_12 = 12;
  localparam th_blink_13 = 13;
  localparam th_blink_14 = 14;
  localparam th_blink_15 = 15;
  localparam th_blink_16 = 16;
  localparam th_blink_17 = 17;
  localparam th_blink_18 = 18;
  localparam th_blink_19 = 19;
  localparam th_blink_20 = 20;
  localparam th_blink_21 = 21;
  localparam th_blink_22 = 22;

  always @(posedge CLK) begin
    if(RST) begin
      th_blink <= th_blink_init;
      done <= 0;
      _th_blink_polarity_259 <= 0;
      _th_blink_tid_260 <= 0;
      _th_myfunc_start[_th_blink_tid_260] <= (0 >> _th_blink_tid_260) & 1'd1;
    end else begin
      case(th_blink)
        th_blink_init: begin
          th_blink <= th_blink_1;
        end
        th_blink_1: begin
          th_blink <= th_blink_2;
        end
        th_blink_2: begin
          if(1) begin
            th_blink <= th_blink_3;
          end else begin
            th_blink <= th_blink_22;
          end
        end
        th_blink_3: begin
          done <= 0;
          th_blink <= th_blink_4;
        end
        th_blink_4: begin
          _th_blink_polarity_259 <= 0;
          th_blink <= th_blink_5;
        end
        th_blink_5: begin
          if(btnC != _th_blink_polarity_259) begin
            th_blink <= th_blink_6;
          end else begin
            th_blink <= th_blink_7;
          end
        end
        th_blink_6: begin
          th_blink <= th_blink_5;
        end
        th_blink_7: begin
          _th_blink_tid_260 <= 0;
          th_blink <= th_blink_8;
        end
        th_blink_8: begin
          if(_th_blink_tid_260 < 64) begin
            th_blink <= th_blink_9;
          end else begin
            th_blink <= th_blink_13;
          end
        end
        th_blink_9: begin
          _th_myfunc_start[_th_blink_tid_260] <= 1;
          th_blink <= th_blink_10;
        end
        th_blink_10: begin
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
        end
        th_blink_11: begin
          _th_myfunc_start[_th_blink_tid_260] <= 0;
          th_blink <= th_blink_12;
        end
        th_blink_12: begin
          _th_blink_tid_260 <= _th_blink_tid_260 + 1;
          th_blink <= th_blink_8;
        end
        th_blink_13: begin
          _th_blink_tid_260 <= 0;
          th_blink <= th_blink_14;
        end
        th_blink_14: begin
          if(_th_blink_tid_260 < 64) begin
            th_blink <= th_blink_15;
          end else begin
            th_blink <= th_blink_17;
          end
        end
        th_blink_15: begin
          if((_th_blink_tid_260 == 0)? th_myfunc_0 == 13 : 
          (_th_blink_tid_260 == 1)? th_myfunc_1 == 13 : 
          (_th_blink_tid_260 == 2)? th_myfunc_2 == 13 : 
          (_th_blink_tid_260 == 3)? th_myfunc_3 == 13 : 
          (_th_blink_tid_260 == 4)? th_myfunc_4 == 13 : 
          (_th_blink_tid_260 == 5)? th_myfunc_5 == 13 : 
          (_th_blink_tid_260 == 6)? th_myfunc_6 == 13 : 
          (_th_blink_tid_260 == 7)? th_myfunc_7 == 13 : 
          (_th_blink_tid_260 == 8)? th_myfunc_8 == 13 : 
          (_th_blink_tid_260 == 9)? th_myfunc_9 == 13 : 
          (_th_blink_tid_260 == 10)? th_myfunc_10 == 13 : 
          (_th_blink_tid_260 == 11)? th_myfunc_11 == 13 : 
          (_th_blink_tid_260 == 12)? th_myfunc_12 == 13 : 
          (_th_blink_tid_260 == 13)? th_myfunc_13 == 13 : 
          (_th_blink_tid_260 == 14)? th_myfunc_14 == 13 : 
          (_th_blink_tid_260 == 15)? th_myfunc_15 == 13 : 
          (_th_blink_tid_260 == 16)? th_myfunc_16 == 13 : 
          (_th_blink_tid_260 == 17)? th_myfunc_17 == 13 : 
          (_th_blink_tid_260 == 18)? th_myfunc_18 == 13 : 
          (_th_blink_tid_260 == 19)? th_myfunc_19 == 13 : 
          (_th_blink_tid_260 == 20)? th_myfunc_20 == 13 : 
          (_th_blink_tid_260 == 21)? th_myfunc_21 == 13 : 
          (_th_blink_tid_260 == 22)? th_myfunc_22 == 13 : 
          (_th_blink_tid_260 == 23)? th_myfunc_23 == 13 : 
          (_th_blink_tid_260 == 24)? th_myfunc_24 == 13 : 
          (_th_blink_tid_260 == 25)? th_myfunc_25 == 13 : 
          (_th_blink_tid_260 == 26)? th_myfunc_26 == 13 : 
          (_th_blink_tid_260 == 27)? th_myfunc_27 == 13 : 
          (_th_blink_tid_260 == 28)? th_myfunc_28 == 13 : 
          (_th_blink_tid_260 == 29)? th_myfunc_29 == 13 : 
          (_th_blink_tid_260 == 30)? th_myfunc_30 == 13 : 
          (_th_blink_tid_260 == 31)? th_myfunc_31 == 13 : 
          (_th_blink_tid_260 == 32)? th_myfunc_32 == 13 : 
          (_th_blink_tid_260 == 33)? th_myfunc_33 == 13 : 
          (_th_blink_tid_260 == 34)? th_myfunc_34 == 13 : 
          (_th_blink_tid_260 == 35)? th_myfunc_35 == 13 : 
          (_th_blink_tid_260 == 36)? th_myfunc_36 == 13 : 
          (_th_blink_tid_260 == 37)? th_myfunc_37 == 13 : 
          (_th_blink_tid_260 == 38)? th_myfunc_38 == 13 : 
          (_th_blink_tid_260 == 39)? th_myfunc_39 == 13 : 
          (_th_blink_tid_260 == 40)? th_myfunc_40 == 13 : 
          (_th_blink_tid_260 == 41)? th_myfunc_41 == 13 : 
          (_th_blink_tid_260 == 42)? th_myfunc_42 == 13 : 
          (_th_blink_tid_260 == 43)? th_myfunc_43 == 13 : 
          (_th_blink_tid_260 == 44)? th_myfunc_44 == 13 : 
          (_th_blink_tid_260 == 45)? th_myfunc_45 == 13 : 
          (_th_blink_tid_260 == 46)? th_myfunc_46 == 13 : 
          (_th_blink_tid_260 == 47)? th_myfunc_47 == 13 : 
          (_th_blink_tid_260 == 48)? th_myfunc_48 == 13 : 
          (_th_blink_tid_260 == 49)? th_myfunc_49 == 13 : 
          (_th_blink_tid_260 == 50)? th_myfunc_50 == 13 : 
          (_th_blink_tid_260 == 51)? th_myfunc_51 == 13 : 
          (_th_blink_tid_260 == 52)? th_myfunc_52 == 13 : 
          (_th_blink_tid_260 == 53)? th_myfunc_53 == 13 : 
          (_th_blink_tid_260 == 54)? th_myfunc_54 == 13 : 
          (_th_blink_tid_260 == 55)? th_myfunc_55 == 13 : 
          (_th_blink_tid_260 == 56)? th_myfunc_56 == 13 : 
          (_th_blink_tid_260 == 57)? th_myfunc_57 == 13 : 
          (_th_blink_tid_260 == 58)? th_myfunc_58 == 13 : 
          (_th_blink_tid_260 == 59)? th_myfunc_59 == 13 : 
          (_th_blink_tid_260 == 60)? th_myfunc_60 == 13 : 
          (_th_blink_tid_260 == 61)? th_myfunc_61 == 13 : 
          (_th_blink_tid_260 == 62)? th_myfunc_62 == 13 : 
          (_th_blink_tid_260 == 63)? th_myfunc_63 == 13 : 0) begin
            th_blink <= th_blink_16;
          end 
        end
        th_blink_16: begin
          _th_blink_tid_260 <= _th_blink_tid_260 + 1;
          th_blink <= th_blink_14;
        end
        th_blink_17: begin
          _th_blink_tid_260 <= 0;
          th_blink <= th_blink_18;
        end
        th_blink_18: begin
          if(_th_blink_tid_260 < 64) begin
            th_blink <= th_blink_19;
          end else begin
            th_blink <= th_blink_20;
          end
        end
        th_blink_19: begin
          _th_blink_tid_260 <= _th_blink_tid_260 + 1;
          th_blink <= th_blink_18;
        end
        th_blink_20: begin
          done <= 1;
          th_blink <= th_blink_21;
        end
        th_blink_21: begin
          th_blink <= th_blink_2;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count <= 0;
    end else begin
      if(th_blink == 1) begin
        count <= 0;
      end 
      if(th_myfunc_0 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_1 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_2 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_3 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_4 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_5 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_6 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_7 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_8 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_9 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_10 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_11 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_12 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_13 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_14 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_15 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_16 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_17 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_18 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_19 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_20 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_21 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_22 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_23 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_24 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_25 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_26 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_27 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_28 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_29 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_30 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_31 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_32 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_33 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_34 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_35 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_36 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_37 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_38 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_39 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_40 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_41 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_42 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_43 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_44 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_45 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_46 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_47 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_48 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_49 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_50 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_51 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_52 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_53 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_54 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_55 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_56 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_57 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_58 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_59 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_60 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_61 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_62 == 9) begin
        count <= count + 1;
      end 
      if(th_myfunc_63 == 9) begin
        count <= count + 1;
      end 
    end
  end

  localparam th_myfunc_0_1 = 1;
  localparam th_myfunc_0_2 = 2;
  localparam th_myfunc_0_3 = 3;
  localparam th_myfunc_0_4 = 4;
  localparam th_myfunc_0_5 = 5;
  localparam th_myfunc_0_6 = 6;
  localparam th_myfunc_0_7 = 7;
  localparam th_myfunc_0_8 = 8;
  localparam th_myfunc_0_9 = 9;
  localparam th_myfunc_0_10 = 10;
  localparam th_myfunc_0_11 = 11;
  localparam th_myfunc_0_12 = 12;
  localparam th_myfunc_0_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_0 <= th_myfunc_0_init;
      _th_myfunc_0_called <= 0;
      _th_myfunc_0_tid_261 <= 0;
      _th_myfunc_0_tid_262 <= 0;
      _th_myfunc_0_time_263 <= 0;
      _th_myfunc_0_i_264 <= 0;
    end else begin
      case(th_myfunc_0)
        th_myfunc_0_init: begin
          if(_th_myfunc_start[0] && (th_blink == 10)) begin
            _th_myfunc_0_called <= 1;
          end 
          if(_th_myfunc_start[0] && (th_blink == 10)) begin
            _th_myfunc_0_tid_261 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[0]) begin
            th_myfunc_0 <= th_myfunc_0_1;
          end 
        end
        th_myfunc_0_1: begin
          _th_myfunc_0_tid_262 <= _th_myfunc_0_tid_261;
          th_myfunc_0 <= th_myfunc_0_2;
        end
        th_myfunc_0_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 0)) begin
            th_myfunc_0 <= th_myfunc_0_3;
          end 
        end
        th_myfunc_0_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 0))) begin
            th_myfunc_0 <= th_myfunc_0_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 0)) begin
            th_myfunc_0 <= th_myfunc_0_4;
          end 
        end
        th_myfunc_0_4: begin
          $display("Thread %d Lock", _th_myfunc_0_tid_262);
          th_myfunc_0 <= th_myfunc_0_5;
        end
        th_myfunc_0_5: begin
          _th_myfunc_0_time_263 <= sw;
          th_myfunc_0 <= th_myfunc_0_6;
        end
        th_myfunc_0_6: begin
          _th_myfunc_0_i_264 <= 0;
          th_myfunc_0 <= th_myfunc_0_7;
        end
        th_myfunc_0_7: begin
          if(_th_myfunc_0_i_264 < _th_myfunc_0_time_263) begin
            th_myfunc_0 <= th_myfunc_0_8;
          end else begin
            th_myfunc_0 <= th_myfunc_0_9;
          end
        end
        th_myfunc_0_8: begin
          _th_myfunc_0_i_264 <= _th_myfunc_0_i_264 + 1;
          th_myfunc_0 <= th_myfunc_0_7;
        end
        th_myfunc_0_9: begin
          th_myfunc_0 <= th_myfunc_0_10;
        end
        th_myfunc_0_10: begin
          $display("Thread %d count = %d", _th_myfunc_0_tid_262, count);
          th_myfunc_0 <= th_myfunc_0_11;
        end
        th_myfunc_0_11: begin
          th_myfunc_0 <= th_myfunc_0_12;
        end
        th_myfunc_0_12: begin
          $display("Thread %d Unlock", _th_myfunc_0_tid_262);
          th_myfunc_0 <= th_myfunc_0_13;
        end
        th_myfunc_0_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 0)) begin
            _th_myfunc_0_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 0)) begin
            th_myfunc_0 <= th_myfunc_0_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_1_1 = 1;
  localparam th_myfunc_1_2 = 2;
  localparam th_myfunc_1_3 = 3;
  localparam th_myfunc_1_4 = 4;
  localparam th_myfunc_1_5 = 5;
  localparam th_myfunc_1_6 = 6;
  localparam th_myfunc_1_7 = 7;
  localparam th_myfunc_1_8 = 8;
  localparam th_myfunc_1_9 = 9;
  localparam th_myfunc_1_10 = 10;
  localparam th_myfunc_1_11 = 11;
  localparam th_myfunc_1_12 = 12;
  localparam th_myfunc_1_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_1 <= th_myfunc_1_init;
      _th_myfunc_1_called <= 0;
      _th_myfunc_1_tid_265 <= 0;
      _th_myfunc_1_tid_266 <= 0;
      _th_myfunc_1_time_267 <= 0;
      _th_myfunc_1_i_268 <= 0;
    end else begin
      case(th_myfunc_1)
        th_myfunc_1_init: begin
          if(_th_myfunc_start[1] && (th_blink == 10)) begin
            _th_myfunc_1_called <= 1;
          end 
          if(_th_myfunc_start[1] && (th_blink == 10)) begin
            _th_myfunc_1_tid_265 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[1]) begin
            th_myfunc_1 <= th_myfunc_1_1;
          end 
        end
        th_myfunc_1_1: begin
          _th_myfunc_1_tid_266 <= _th_myfunc_1_tid_265;
          th_myfunc_1 <= th_myfunc_1_2;
        end
        th_myfunc_1_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 1)) begin
            th_myfunc_1 <= th_myfunc_1_3;
          end 
        end
        th_myfunc_1_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 1))) begin
            th_myfunc_1 <= th_myfunc_1_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 1)) begin
            th_myfunc_1 <= th_myfunc_1_4;
          end 
        end
        th_myfunc_1_4: begin
          $display("Thread %d Lock", _th_myfunc_1_tid_266);
          th_myfunc_1 <= th_myfunc_1_5;
        end
        th_myfunc_1_5: begin
          _th_myfunc_1_time_267 <= sw;
          th_myfunc_1 <= th_myfunc_1_6;
        end
        th_myfunc_1_6: begin
          _th_myfunc_1_i_268 <= 0;
          th_myfunc_1 <= th_myfunc_1_7;
        end
        th_myfunc_1_7: begin
          if(_th_myfunc_1_i_268 < _th_myfunc_1_time_267) begin
            th_myfunc_1 <= th_myfunc_1_8;
          end else begin
            th_myfunc_1 <= th_myfunc_1_9;
          end
        end
        th_myfunc_1_8: begin
          _th_myfunc_1_i_268 <= _th_myfunc_1_i_268 + 1;
          th_myfunc_1 <= th_myfunc_1_7;
        end
        th_myfunc_1_9: begin
          th_myfunc_1 <= th_myfunc_1_10;
        end
        th_myfunc_1_10: begin
          $display("Thread %d count = %d", _th_myfunc_1_tid_266, count);
          th_myfunc_1 <= th_myfunc_1_11;
        end
        th_myfunc_1_11: begin
          th_myfunc_1 <= th_myfunc_1_12;
        end
        th_myfunc_1_12: begin
          $display("Thread %d Unlock", _th_myfunc_1_tid_266);
          th_myfunc_1 <= th_myfunc_1_13;
        end
        th_myfunc_1_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 1)) begin
            _th_myfunc_1_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 1)) begin
            th_myfunc_1 <= th_myfunc_1_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_2_1 = 1;
  localparam th_myfunc_2_2 = 2;
  localparam th_myfunc_2_3 = 3;
  localparam th_myfunc_2_4 = 4;
  localparam th_myfunc_2_5 = 5;
  localparam th_myfunc_2_6 = 6;
  localparam th_myfunc_2_7 = 7;
  localparam th_myfunc_2_8 = 8;
  localparam th_myfunc_2_9 = 9;
  localparam th_myfunc_2_10 = 10;
  localparam th_myfunc_2_11 = 11;
  localparam th_myfunc_2_12 = 12;
  localparam th_myfunc_2_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_2 <= th_myfunc_2_init;
      _th_myfunc_2_called <= 0;
      _th_myfunc_2_tid_269 <= 0;
      _th_myfunc_2_tid_270 <= 0;
      _th_myfunc_2_time_271 <= 0;
      _th_myfunc_2_i_272 <= 0;
    end else begin
      case(th_myfunc_2)
        th_myfunc_2_init: begin
          if(_th_myfunc_start[2] && (th_blink == 10)) begin
            _th_myfunc_2_called <= 1;
          end 
          if(_th_myfunc_start[2] && (th_blink == 10)) begin
            _th_myfunc_2_tid_269 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[2]) begin
            th_myfunc_2 <= th_myfunc_2_1;
          end 
        end
        th_myfunc_2_1: begin
          _th_myfunc_2_tid_270 <= _th_myfunc_2_tid_269;
          th_myfunc_2 <= th_myfunc_2_2;
        end
        th_myfunc_2_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 2)) begin
            th_myfunc_2 <= th_myfunc_2_3;
          end 
        end
        th_myfunc_2_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 2))) begin
            th_myfunc_2 <= th_myfunc_2_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 2)) begin
            th_myfunc_2 <= th_myfunc_2_4;
          end 
        end
        th_myfunc_2_4: begin
          $display("Thread %d Lock", _th_myfunc_2_tid_270);
          th_myfunc_2 <= th_myfunc_2_5;
        end
        th_myfunc_2_5: begin
          _th_myfunc_2_time_271 <= sw;
          th_myfunc_2 <= th_myfunc_2_6;
        end
        th_myfunc_2_6: begin
          _th_myfunc_2_i_272 <= 0;
          th_myfunc_2 <= th_myfunc_2_7;
        end
        th_myfunc_2_7: begin
          if(_th_myfunc_2_i_272 < _th_myfunc_2_time_271) begin
            th_myfunc_2 <= th_myfunc_2_8;
          end else begin
            th_myfunc_2 <= th_myfunc_2_9;
          end
        end
        th_myfunc_2_8: begin
          _th_myfunc_2_i_272 <= _th_myfunc_2_i_272 + 1;
          th_myfunc_2 <= th_myfunc_2_7;
        end
        th_myfunc_2_9: begin
          th_myfunc_2 <= th_myfunc_2_10;
        end
        th_myfunc_2_10: begin
          $display("Thread %d count = %d", _th_myfunc_2_tid_270, count);
          th_myfunc_2 <= th_myfunc_2_11;
        end
        th_myfunc_2_11: begin
          th_myfunc_2 <= th_myfunc_2_12;
        end
        th_myfunc_2_12: begin
          $display("Thread %d Unlock", _th_myfunc_2_tid_270);
          th_myfunc_2 <= th_myfunc_2_13;
        end
        th_myfunc_2_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 2)) begin
            _th_myfunc_2_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 2)) begin
            th_myfunc_2 <= th_myfunc_2_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_3_1 = 1;
  localparam th_myfunc_3_2 = 2;
  localparam th_myfunc_3_3 = 3;
  localparam th_myfunc_3_4 = 4;
  localparam th_myfunc_3_5 = 5;
  localparam th_myfunc_3_6 = 6;
  localparam th_myfunc_3_7 = 7;
  localparam th_myfunc_3_8 = 8;
  localparam th_myfunc_3_9 = 9;
  localparam th_myfunc_3_10 = 10;
  localparam th_myfunc_3_11 = 11;
  localparam th_myfunc_3_12 = 12;
  localparam th_myfunc_3_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_3 <= th_myfunc_3_init;
      _th_myfunc_3_called <= 0;
      _th_myfunc_3_tid_273 <= 0;
      _th_myfunc_3_tid_274 <= 0;
      _th_myfunc_3_time_275 <= 0;
      _th_myfunc_3_i_276 <= 0;
    end else begin
      case(th_myfunc_3)
        th_myfunc_3_init: begin
          if(_th_myfunc_start[3] && (th_blink == 10)) begin
            _th_myfunc_3_called <= 1;
          end 
          if(_th_myfunc_start[3] && (th_blink == 10)) begin
            _th_myfunc_3_tid_273 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[3]) begin
            th_myfunc_3 <= th_myfunc_3_1;
          end 
        end
        th_myfunc_3_1: begin
          _th_myfunc_3_tid_274 <= _th_myfunc_3_tid_273;
          th_myfunc_3 <= th_myfunc_3_2;
        end
        th_myfunc_3_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 3)) begin
            th_myfunc_3 <= th_myfunc_3_3;
          end 
        end
        th_myfunc_3_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 3))) begin
            th_myfunc_3 <= th_myfunc_3_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 3)) begin
            th_myfunc_3 <= th_myfunc_3_4;
          end 
        end
        th_myfunc_3_4: begin
          $display("Thread %d Lock", _th_myfunc_3_tid_274);
          th_myfunc_3 <= th_myfunc_3_5;
        end
        th_myfunc_3_5: begin
          _th_myfunc_3_time_275 <= sw;
          th_myfunc_3 <= th_myfunc_3_6;
        end
        th_myfunc_3_6: begin
          _th_myfunc_3_i_276 <= 0;
          th_myfunc_3 <= th_myfunc_3_7;
        end
        th_myfunc_3_7: begin
          if(_th_myfunc_3_i_276 < _th_myfunc_3_time_275) begin
            th_myfunc_3 <= th_myfunc_3_8;
          end else begin
            th_myfunc_3 <= th_myfunc_3_9;
          end
        end
        th_myfunc_3_8: begin
          _th_myfunc_3_i_276 <= _th_myfunc_3_i_276 + 1;
          th_myfunc_3 <= th_myfunc_3_7;
        end
        th_myfunc_3_9: begin
          th_myfunc_3 <= th_myfunc_3_10;
        end
        th_myfunc_3_10: begin
          $display("Thread %d count = %d", _th_myfunc_3_tid_274, count);
          th_myfunc_3 <= th_myfunc_3_11;
        end
        th_myfunc_3_11: begin
          th_myfunc_3 <= th_myfunc_3_12;
        end
        th_myfunc_3_12: begin
          $display("Thread %d Unlock", _th_myfunc_3_tid_274);
          th_myfunc_3 <= th_myfunc_3_13;
        end
        th_myfunc_3_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 3)) begin
            _th_myfunc_3_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 3)) begin
            th_myfunc_3 <= th_myfunc_3_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_4_1 = 1;
  localparam th_myfunc_4_2 = 2;
  localparam th_myfunc_4_3 = 3;
  localparam th_myfunc_4_4 = 4;
  localparam th_myfunc_4_5 = 5;
  localparam th_myfunc_4_6 = 6;
  localparam th_myfunc_4_7 = 7;
  localparam th_myfunc_4_8 = 8;
  localparam th_myfunc_4_9 = 9;
  localparam th_myfunc_4_10 = 10;
  localparam th_myfunc_4_11 = 11;
  localparam th_myfunc_4_12 = 12;
  localparam th_myfunc_4_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_4 <= th_myfunc_4_init;
      _th_myfunc_4_called <= 0;
      _th_myfunc_4_tid_277 <= 0;
      _th_myfunc_4_tid_278 <= 0;
      _th_myfunc_4_time_279 <= 0;
      _th_myfunc_4_i_280 <= 0;
    end else begin
      case(th_myfunc_4)
        th_myfunc_4_init: begin
          if(_th_myfunc_start[4] && (th_blink == 10)) begin
            _th_myfunc_4_called <= 1;
          end 
          if(_th_myfunc_start[4] && (th_blink == 10)) begin
            _th_myfunc_4_tid_277 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[4]) begin
            th_myfunc_4 <= th_myfunc_4_1;
          end 
        end
        th_myfunc_4_1: begin
          _th_myfunc_4_tid_278 <= _th_myfunc_4_tid_277;
          th_myfunc_4 <= th_myfunc_4_2;
        end
        th_myfunc_4_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 4)) begin
            th_myfunc_4 <= th_myfunc_4_3;
          end 
        end
        th_myfunc_4_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 4))) begin
            th_myfunc_4 <= th_myfunc_4_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 4)) begin
            th_myfunc_4 <= th_myfunc_4_4;
          end 
        end
        th_myfunc_4_4: begin
          $display("Thread %d Lock", _th_myfunc_4_tid_278);
          th_myfunc_4 <= th_myfunc_4_5;
        end
        th_myfunc_4_5: begin
          _th_myfunc_4_time_279 <= sw;
          th_myfunc_4 <= th_myfunc_4_6;
        end
        th_myfunc_4_6: begin
          _th_myfunc_4_i_280 <= 0;
          th_myfunc_4 <= th_myfunc_4_7;
        end
        th_myfunc_4_7: begin
          if(_th_myfunc_4_i_280 < _th_myfunc_4_time_279) begin
            th_myfunc_4 <= th_myfunc_4_8;
          end else begin
            th_myfunc_4 <= th_myfunc_4_9;
          end
        end
        th_myfunc_4_8: begin
          _th_myfunc_4_i_280 <= _th_myfunc_4_i_280 + 1;
          th_myfunc_4 <= th_myfunc_4_7;
        end
        th_myfunc_4_9: begin
          th_myfunc_4 <= th_myfunc_4_10;
        end
        th_myfunc_4_10: begin
          $display("Thread %d count = %d", _th_myfunc_4_tid_278, count);
          th_myfunc_4 <= th_myfunc_4_11;
        end
        th_myfunc_4_11: begin
          th_myfunc_4 <= th_myfunc_4_12;
        end
        th_myfunc_4_12: begin
          $display("Thread %d Unlock", _th_myfunc_4_tid_278);
          th_myfunc_4 <= th_myfunc_4_13;
        end
        th_myfunc_4_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 4)) begin
            _th_myfunc_4_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 4)) begin
            th_myfunc_4 <= th_myfunc_4_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_5_1 = 1;
  localparam th_myfunc_5_2 = 2;
  localparam th_myfunc_5_3 = 3;
  localparam th_myfunc_5_4 = 4;
  localparam th_myfunc_5_5 = 5;
  localparam th_myfunc_5_6 = 6;
  localparam th_myfunc_5_7 = 7;
  localparam th_myfunc_5_8 = 8;
  localparam th_myfunc_5_9 = 9;
  localparam th_myfunc_5_10 = 10;
  localparam th_myfunc_5_11 = 11;
  localparam th_myfunc_5_12 = 12;
  localparam th_myfunc_5_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_5 <= th_myfunc_5_init;
      _th_myfunc_5_called <= 0;
      _th_myfunc_5_tid_281 <= 0;
      _th_myfunc_5_tid_282 <= 0;
      _th_myfunc_5_time_283 <= 0;
      _th_myfunc_5_i_284 <= 0;
    end else begin
      case(th_myfunc_5)
        th_myfunc_5_init: begin
          if(_th_myfunc_start[5] && (th_blink == 10)) begin
            _th_myfunc_5_called <= 1;
          end 
          if(_th_myfunc_start[5] && (th_blink == 10)) begin
            _th_myfunc_5_tid_281 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[5]) begin
            th_myfunc_5 <= th_myfunc_5_1;
          end 
        end
        th_myfunc_5_1: begin
          _th_myfunc_5_tid_282 <= _th_myfunc_5_tid_281;
          th_myfunc_5 <= th_myfunc_5_2;
        end
        th_myfunc_5_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 5)) begin
            th_myfunc_5 <= th_myfunc_5_3;
          end 
        end
        th_myfunc_5_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 5))) begin
            th_myfunc_5 <= th_myfunc_5_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 5)) begin
            th_myfunc_5 <= th_myfunc_5_4;
          end 
        end
        th_myfunc_5_4: begin
          $display("Thread %d Lock", _th_myfunc_5_tid_282);
          th_myfunc_5 <= th_myfunc_5_5;
        end
        th_myfunc_5_5: begin
          _th_myfunc_5_time_283 <= sw;
          th_myfunc_5 <= th_myfunc_5_6;
        end
        th_myfunc_5_6: begin
          _th_myfunc_5_i_284 <= 0;
          th_myfunc_5 <= th_myfunc_5_7;
        end
        th_myfunc_5_7: begin
          if(_th_myfunc_5_i_284 < _th_myfunc_5_time_283) begin
            th_myfunc_5 <= th_myfunc_5_8;
          end else begin
            th_myfunc_5 <= th_myfunc_5_9;
          end
        end
        th_myfunc_5_8: begin
          _th_myfunc_5_i_284 <= _th_myfunc_5_i_284 + 1;
          th_myfunc_5 <= th_myfunc_5_7;
        end
        th_myfunc_5_9: begin
          th_myfunc_5 <= th_myfunc_5_10;
        end
        th_myfunc_5_10: begin
          $display("Thread %d count = %d", _th_myfunc_5_tid_282, count);
          th_myfunc_5 <= th_myfunc_5_11;
        end
        th_myfunc_5_11: begin
          th_myfunc_5 <= th_myfunc_5_12;
        end
        th_myfunc_5_12: begin
          $display("Thread %d Unlock", _th_myfunc_5_tid_282);
          th_myfunc_5 <= th_myfunc_5_13;
        end
        th_myfunc_5_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 5)) begin
            _th_myfunc_5_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 5)) begin
            th_myfunc_5 <= th_myfunc_5_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_6_1 = 1;
  localparam th_myfunc_6_2 = 2;
  localparam th_myfunc_6_3 = 3;
  localparam th_myfunc_6_4 = 4;
  localparam th_myfunc_6_5 = 5;
  localparam th_myfunc_6_6 = 6;
  localparam th_myfunc_6_7 = 7;
  localparam th_myfunc_6_8 = 8;
  localparam th_myfunc_6_9 = 9;
  localparam th_myfunc_6_10 = 10;
  localparam th_myfunc_6_11 = 11;
  localparam th_myfunc_6_12 = 12;
  localparam th_myfunc_6_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_6 <= th_myfunc_6_init;
      _th_myfunc_6_called <= 0;
      _th_myfunc_6_tid_285 <= 0;
      _th_myfunc_6_tid_286 <= 0;
      _th_myfunc_6_time_287 <= 0;
      _th_myfunc_6_i_288 <= 0;
    end else begin
      case(th_myfunc_6)
        th_myfunc_6_init: begin
          if(_th_myfunc_start[6] && (th_blink == 10)) begin
            _th_myfunc_6_called <= 1;
          end 
          if(_th_myfunc_start[6] && (th_blink == 10)) begin
            _th_myfunc_6_tid_285 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[6]) begin
            th_myfunc_6 <= th_myfunc_6_1;
          end 
        end
        th_myfunc_6_1: begin
          _th_myfunc_6_tid_286 <= _th_myfunc_6_tid_285;
          th_myfunc_6 <= th_myfunc_6_2;
        end
        th_myfunc_6_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 6)) begin
            th_myfunc_6 <= th_myfunc_6_3;
          end 
        end
        th_myfunc_6_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 6))) begin
            th_myfunc_6 <= th_myfunc_6_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 6)) begin
            th_myfunc_6 <= th_myfunc_6_4;
          end 
        end
        th_myfunc_6_4: begin
          $display("Thread %d Lock", _th_myfunc_6_tid_286);
          th_myfunc_6 <= th_myfunc_6_5;
        end
        th_myfunc_6_5: begin
          _th_myfunc_6_time_287 <= sw;
          th_myfunc_6 <= th_myfunc_6_6;
        end
        th_myfunc_6_6: begin
          _th_myfunc_6_i_288 <= 0;
          th_myfunc_6 <= th_myfunc_6_7;
        end
        th_myfunc_6_7: begin
          if(_th_myfunc_6_i_288 < _th_myfunc_6_time_287) begin
            th_myfunc_6 <= th_myfunc_6_8;
          end else begin
            th_myfunc_6 <= th_myfunc_6_9;
          end
        end
        th_myfunc_6_8: begin
          _th_myfunc_6_i_288 <= _th_myfunc_6_i_288 + 1;
          th_myfunc_6 <= th_myfunc_6_7;
        end
        th_myfunc_6_9: begin
          th_myfunc_6 <= th_myfunc_6_10;
        end
        th_myfunc_6_10: begin
          $display("Thread %d count = %d", _th_myfunc_6_tid_286, count);
          th_myfunc_6 <= th_myfunc_6_11;
        end
        th_myfunc_6_11: begin
          th_myfunc_6 <= th_myfunc_6_12;
        end
        th_myfunc_6_12: begin
          $display("Thread %d Unlock", _th_myfunc_6_tid_286);
          th_myfunc_6 <= th_myfunc_6_13;
        end
        th_myfunc_6_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 6)) begin
            _th_myfunc_6_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 6)) begin
            th_myfunc_6 <= th_myfunc_6_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_7_1 = 1;
  localparam th_myfunc_7_2 = 2;
  localparam th_myfunc_7_3 = 3;
  localparam th_myfunc_7_4 = 4;
  localparam th_myfunc_7_5 = 5;
  localparam th_myfunc_7_6 = 6;
  localparam th_myfunc_7_7 = 7;
  localparam th_myfunc_7_8 = 8;
  localparam th_myfunc_7_9 = 9;
  localparam th_myfunc_7_10 = 10;
  localparam th_myfunc_7_11 = 11;
  localparam th_myfunc_7_12 = 12;
  localparam th_myfunc_7_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_7 <= th_myfunc_7_init;
      _th_myfunc_7_called <= 0;
      _th_myfunc_7_tid_289 <= 0;
      _th_myfunc_7_tid_290 <= 0;
      _th_myfunc_7_time_291 <= 0;
      _th_myfunc_7_i_292 <= 0;
    end else begin
      case(th_myfunc_7)
        th_myfunc_7_init: begin
          if(_th_myfunc_start[7] && (th_blink == 10)) begin
            _th_myfunc_7_called <= 1;
          end 
          if(_th_myfunc_start[7] && (th_blink == 10)) begin
            _th_myfunc_7_tid_289 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[7]) begin
            th_myfunc_7 <= th_myfunc_7_1;
          end 
        end
        th_myfunc_7_1: begin
          _th_myfunc_7_tid_290 <= _th_myfunc_7_tid_289;
          th_myfunc_7 <= th_myfunc_7_2;
        end
        th_myfunc_7_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 7)) begin
            th_myfunc_7 <= th_myfunc_7_3;
          end 
        end
        th_myfunc_7_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 7))) begin
            th_myfunc_7 <= th_myfunc_7_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 7)) begin
            th_myfunc_7 <= th_myfunc_7_4;
          end 
        end
        th_myfunc_7_4: begin
          $display("Thread %d Lock", _th_myfunc_7_tid_290);
          th_myfunc_7 <= th_myfunc_7_5;
        end
        th_myfunc_7_5: begin
          _th_myfunc_7_time_291 <= sw;
          th_myfunc_7 <= th_myfunc_7_6;
        end
        th_myfunc_7_6: begin
          _th_myfunc_7_i_292 <= 0;
          th_myfunc_7 <= th_myfunc_7_7;
        end
        th_myfunc_7_7: begin
          if(_th_myfunc_7_i_292 < _th_myfunc_7_time_291) begin
            th_myfunc_7 <= th_myfunc_7_8;
          end else begin
            th_myfunc_7 <= th_myfunc_7_9;
          end
        end
        th_myfunc_7_8: begin
          _th_myfunc_7_i_292 <= _th_myfunc_7_i_292 + 1;
          th_myfunc_7 <= th_myfunc_7_7;
        end
        th_myfunc_7_9: begin
          th_myfunc_7 <= th_myfunc_7_10;
        end
        th_myfunc_7_10: begin
          $display("Thread %d count = %d", _th_myfunc_7_tid_290, count);
          th_myfunc_7 <= th_myfunc_7_11;
        end
        th_myfunc_7_11: begin
          th_myfunc_7 <= th_myfunc_7_12;
        end
        th_myfunc_7_12: begin
          $display("Thread %d Unlock", _th_myfunc_7_tid_290);
          th_myfunc_7 <= th_myfunc_7_13;
        end
        th_myfunc_7_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 7)) begin
            _th_myfunc_7_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 7)) begin
            th_myfunc_7 <= th_myfunc_7_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_8_1 = 1;
  localparam th_myfunc_8_2 = 2;
  localparam th_myfunc_8_3 = 3;
  localparam th_myfunc_8_4 = 4;
  localparam th_myfunc_8_5 = 5;
  localparam th_myfunc_8_6 = 6;
  localparam th_myfunc_8_7 = 7;
  localparam th_myfunc_8_8 = 8;
  localparam th_myfunc_8_9 = 9;
  localparam th_myfunc_8_10 = 10;
  localparam th_myfunc_8_11 = 11;
  localparam th_myfunc_8_12 = 12;
  localparam th_myfunc_8_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_8 <= th_myfunc_8_init;
      _th_myfunc_8_called <= 0;
      _th_myfunc_8_tid_293 <= 0;
      _th_myfunc_8_tid_294 <= 0;
      _th_myfunc_8_time_295 <= 0;
      _th_myfunc_8_i_296 <= 0;
    end else begin
      case(th_myfunc_8)
        th_myfunc_8_init: begin
          if(_th_myfunc_start[8] && (th_blink == 10)) begin
            _th_myfunc_8_called <= 1;
          end 
          if(_th_myfunc_start[8] && (th_blink == 10)) begin
            _th_myfunc_8_tid_293 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[8]) begin
            th_myfunc_8 <= th_myfunc_8_1;
          end 
        end
        th_myfunc_8_1: begin
          _th_myfunc_8_tid_294 <= _th_myfunc_8_tid_293;
          th_myfunc_8 <= th_myfunc_8_2;
        end
        th_myfunc_8_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 8)) begin
            th_myfunc_8 <= th_myfunc_8_3;
          end 
        end
        th_myfunc_8_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 8))) begin
            th_myfunc_8 <= th_myfunc_8_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 8)) begin
            th_myfunc_8 <= th_myfunc_8_4;
          end 
        end
        th_myfunc_8_4: begin
          $display("Thread %d Lock", _th_myfunc_8_tid_294);
          th_myfunc_8 <= th_myfunc_8_5;
        end
        th_myfunc_8_5: begin
          _th_myfunc_8_time_295 <= sw;
          th_myfunc_8 <= th_myfunc_8_6;
        end
        th_myfunc_8_6: begin
          _th_myfunc_8_i_296 <= 0;
          th_myfunc_8 <= th_myfunc_8_7;
        end
        th_myfunc_8_7: begin
          if(_th_myfunc_8_i_296 < _th_myfunc_8_time_295) begin
            th_myfunc_8 <= th_myfunc_8_8;
          end else begin
            th_myfunc_8 <= th_myfunc_8_9;
          end
        end
        th_myfunc_8_8: begin
          _th_myfunc_8_i_296 <= _th_myfunc_8_i_296 + 1;
          th_myfunc_8 <= th_myfunc_8_7;
        end
        th_myfunc_8_9: begin
          th_myfunc_8 <= th_myfunc_8_10;
        end
        th_myfunc_8_10: begin
          $display("Thread %d count = %d", _th_myfunc_8_tid_294, count);
          th_myfunc_8 <= th_myfunc_8_11;
        end
        th_myfunc_8_11: begin
          th_myfunc_8 <= th_myfunc_8_12;
        end
        th_myfunc_8_12: begin
          $display("Thread %d Unlock", _th_myfunc_8_tid_294);
          th_myfunc_8 <= th_myfunc_8_13;
        end
        th_myfunc_8_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 8)) begin
            _th_myfunc_8_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 8)) begin
            th_myfunc_8 <= th_myfunc_8_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_9_1 = 1;
  localparam th_myfunc_9_2 = 2;
  localparam th_myfunc_9_3 = 3;
  localparam th_myfunc_9_4 = 4;
  localparam th_myfunc_9_5 = 5;
  localparam th_myfunc_9_6 = 6;
  localparam th_myfunc_9_7 = 7;
  localparam th_myfunc_9_8 = 8;
  localparam th_myfunc_9_9 = 9;
  localparam th_myfunc_9_10 = 10;
  localparam th_myfunc_9_11 = 11;
  localparam th_myfunc_9_12 = 12;
  localparam th_myfunc_9_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_9 <= th_myfunc_9_init;
      _th_myfunc_9_called <= 0;
      _th_myfunc_9_tid_297 <= 0;
      _th_myfunc_9_tid_298 <= 0;
      _th_myfunc_9_time_299 <= 0;
      _th_myfunc_9_i_300 <= 0;
    end else begin
      case(th_myfunc_9)
        th_myfunc_9_init: begin
          if(_th_myfunc_start[9] && (th_blink == 10)) begin
            _th_myfunc_9_called <= 1;
          end 
          if(_th_myfunc_start[9] && (th_blink == 10)) begin
            _th_myfunc_9_tid_297 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[9]) begin
            th_myfunc_9 <= th_myfunc_9_1;
          end 
        end
        th_myfunc_9_1: begin
          _th_myfunc_9_tid_298 <= _th_myfunc_9_tid_297;
          th_myfunc_9 <= th_myfunc_9_2;
        end
        th_myfunc_9_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 9)) begin
            th_myfunc_9 <= th_myfunc_9_3;
          end 
        end
        th_myfunc_9_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 9))) begin
            th_myfunc_9 <= th_myfunc_9_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 9)) begin
            th_myfunc_9 <= th_myfunc_9_4;
          end 
        end
        th_myfunc_9_4: begin
          $display("Thread %d Lock", _th_myfunc_9_tid_298);
          th_myfunc_9 <= th_myfunc_9_5;
        end
        th_myfunc_9_5: begin
          _th_myfunc_9_time_299 <= sw;
          th_myfunc_9 <= th_myfunc_9_6;
        end
        th_myfunc_9_6: begin
          _th_myfunc_9_i_300 <= 0;
          th_myfunc_9 <= th_myfunc_9_7;
        end
        th_myfunc_9_7: begin
          if(_th_myfunc_9_i_300 < _th_myfunc_9_time_299) begin
            th_myfunc_9 <= th_myfunc_9_8;
          end else begin
            th_myfunc_9 <= th_myfunc_9_9;
          end
        end
        th_myfunc_9_8: begin
          _th_myfunc_9_i_300 <= _th_myfunc_9_i_300 + 1;
          th_myfunc_9 <= th_myfunc_9_7;
        end
        th_myfunc_9_9: begin
          th_myfunc_9 <= th_myfunc_9_10;
        end
        th_myfunc_9_10: begin
          $display("Thread %d count = %d", _th_myfunc_9_tid_298, count);
          th_myfunc_9 <= th_myfunc_9_11;
        end
        th_myfunc_9_11: begin
          th_myfunc_9 <= th_myfunc_9_12;
        end
        th_myfunc_9_12: begin
          $display("Thread %d Unlock", _th_myfunc_9_tid_298);
          th_myfunc_9 <= th_myfunc_9_13;
        end
        th_myfunc_9_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 9)) begin
            _th_myfunc_9_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 9)) begin
            th_myfunc_9 <= th_myfunc_9_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_10_1 = 1;
  localparam th_myfunc_10_2 = 2;
  localparam th_myfunc_10_3 = 3;
  localparam th_myfunc_10_4 = 4;
  localparam th_myfunc_10_5 = 5;
  localparam th_myfunc_10_6 = 6;
  localparam th_myfunc_10_7 = 7;
  localparam th_myfunc_10_8 = 8;
  localparam th_myfunc_10_9 = 9;
  localparam th_myfunc_10_10 = 10;
  localparam th_myfunc_10_11 = 11;
  localparam th_myfunc_10_12 = 12;
  localparam th_myfunc_10_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_10 <= th_myfunc_10_init;
      _th_myfunc_10_called <= 0;
      _th_myfunc_10_tid_301 <= 0;
      _th_myfunc_10_tid_302 <= 0;
      _th_myfunc_10_time_303 <= 0;
      _th_myfunc_10_i_304 <= 0;
    end else begin
      case(th_myfunc_10)
        th_myfunc_10_init: begin
          if(_th_myfunc_start[10] && (th_blink == 10)) begin
            _th_myfunc_10_called <= 1;
          end 
          if(_th_myfunc_start[10] && (th_blink == 10)) begin
            _th_myfunc_10_tid_301 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[10]) begin
            th_myfunc_10 <= th_myfunc_10_1;
          end 
        end
        th_myfunc_10_1: begin
          _th_myfunc_10_tid_302 <= _th_myfunc_10_tid_301;
          th_myfunc_10 <= th_myfunc_10_2;
        end
        th_myfunc_10_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 10)) begin
            th_myfunc_10 <= th_myfunc_10_3;
          end 
        end
        th_myfunc_10_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 10))) begin
            th_myfunc_10 <= th_myfunc_10_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 10)) begin
            th_myfunc_10 <= th_myfunc_10_4;
          end 
        end
        th_myfunc_10_4: begin
          $display("Thread %d Lock", _th_myfunc_10_tid_302);
          th_myfunc_10 <= th_myfunc_10_5;
        end
        th_myfunc_10_5: begin
          _th_myfunc_10_time_303 <= sw;
          th_myfunc_10 <= th_myfunc_10_6;
        end
        th_myfunc_10_6: begin
          _th_myfunc_10_i_304 <= 0;
          th_myfunc_10 <= th_myfunc_10_7;
        end
        th_myfunc_10_7: begin
          if(_th_myfunc_10_i_304 < _th_myfunc_10_time_303) begin
            th_myfunc_10 <= th_myfunc_10_8;
          end else begin
            th_myfunc_10 <= th_myfunc_10_9;
          end
        end
        th_myfunc_10_8: begin
          _th_myfunc_10_i_304 <= _th_myfunc_10_i_304 + 1;
          th_myfunc_10 <= th_myfunc_10_7;
        end
        th_myfunc_10_9: begin
          th_myfunc_10 <= th_myfunc_10_10;
        end
        th_myfunc_10_10: begin
          $display("Thread %d count = %d", _th_myfunc_10_tid_302, count);
          th_myfunc_10 <= th_myfunc_10_11;
        end
        th_myfunc_10_11: begin
          th_myfunc_10 <= th_myfunc_10_12;
        end
        th_myfunc_10_12: begin
          $display("Thread %d Unlock", _th_myfunc_10_tid_302);
          th_myfunc_10 <= th_myfunc_10_13;
        end
        th_myfunc_10_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 10)) begin
            _th_myfunc_10_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 10)) begin
            th_myfunc_10 <= th_myfunc_10_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_11_1 = 1;
  localparam th_myfunc_11_2 = 2;
  localparam th_myfunc_11_3 = 3;
  localparam th_myfunc_11_4 = 4;
  localparam th_myfunc_11_5 = 5;
  localparam th_myfunc_11_6 = 6;
  localparam th_myfunc_11_7 = 7;
  localparam th_myfunc_11_8 = 8;
  localparam th_myfunc_11_9 = 9;
  localparam th_myfunc_11_10 = 10;
  localparam th_myfunc_11_11 = 11;
  localparam th_myfunc_11_12 = 12;
  localparam th_myfunc_11_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_11 <= th_myfunc_11_init;
      _th_myfunc_11_called <= 0;
      _th_myfunc_11_tid_305 <= 0;
      _th_myfunc_11_tid_306 <= 0;
      _th_myfunc_11_time_307 <= 0;
      _th_myfunc_11_i_308 <= 0;
    end else begin
      case(th_myfunc_11)
        th_myfunc_11_init: begin
          if(_th_myfunc_start[11] && (th_blink == 10)) begin
            _th_myfunc_11_called <= 1;
          end 
          if(_th_myfunc_start[11] && (th_blink == 10)) begin
            _th_myfunc_11_tid_305 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[11]) begin
            th_myfunc_11 <= th_myfunc_11_1;
          end 
        end
        th_myfunc_11_1: begin
          _th_myfunc_11_tid_306 <= _th_myfunc_11_tid_305;
          th_myfunc_11 <= th_myfunc_11_2;
        end
        th_myfunc_11_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 11)) begin
            th_myfunc_11 <= th_myfunc_11_3;
          end 
        end
        th_myfunc_11_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 11))) begin
            th_myfunc_11 <= th_myfunc_11_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 11)) begin
            th_myfunc_11 <= th_myfunc_11_4;
          end 
        end
        th_myfunc_11_4: begin
          $display("Thread %d Lock", _th_myfunc_11_tid_306);
          th_myfunc_11 <= th_myfunc_11_5;
        end
        th_myfunc_11_5: begin
          _th_myfunc_11_time_307 <= sw;
          th_myfunc_11 <= th_myfunc_11_6;
        end
        th_myfunc_11_6: begin
          _th_myfunc_11_i_308 <= 0;
          th_myfunc_11 <= th_myfunc_11_7;
        end
        th_myfunc_11_7: begin
          if(_th_myfunc_11_i_308 < _th_myfunc_11_time_307) begin
            th_myfunc_11 <= th_myfunc_11_8;
          end else begin
            th_myfunc_11 <= th_myfunc_11_9;
          end
        end
        th_myfunc_11_8: begin
          _th_myfunc_11_i_308 <= _th_myfunc_11_i_308 + 1;
          th_myfunc_11 <= th_myfunc_11_7;
        end
        th_myfunc_11_9: begin
          th_myfunc_11 <= th_myfunc_11_10;
        end
        th_myfunc_11_10: begin
          $display("Thread %d count = %d", _th_myfunc_11_tid_306, count);
          th_myfunc_11 <= th_myfunc_11_11;
        end
        th_myfunc_11_11: begin
          th_myfunc_11 <= th_myfunc_11_12;
        end
        th_myfunc_11_12: begin
          $display("Thread %d Unlock", _th_myfunc_11_tid_306);
          th_myfunc_11 <= th_myfunc_11_13;
        end
        th_myfunc_11_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 11)) begin
            _th_myfunc_11_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 11)) begin
            th_myfunc_11 <= th_myfunc_11_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_12_1 = 1;
  localparam th_myfunc_12_2 = 2;
  localparam th_myfunc_12_3 = 3;
  localparam th_myfunc_12_4 = 4;
  localparam th_myfunc_12_5 = 5;
  localparam th_myfunc_12_6 = 6;
  localparam th_myfunc_12_7 = 7;
  localparam th_myfunc_12_8 = 8;
  localparam th_myfunc_12_9 = 9;
  localparam th_myfunc_12_10 = 10;
  localparam th_myfunc_12_11 = 11;
  localparam th_myfunc_12_12 = 12;
  localparam th_myfunc_12_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_12 <= th_myfunc_12_init;
      _th_myfunc_12_called <= 0;
      _th_myfunc_12_tid_309 <= 0;
      _th_myfunc_12_tid_310 <= 0;
      _th_myfunc_12_time_311 <= 0;
      _th_myfunc_12_i_312 <= 0;
    end else begin
      case(th_myfunc_12)
        th_myfunc_12_init: begin
          if(_th_myfunc_start[12] && (th_blink == 10)) begin
            _th_myfunc_12_called <= 1;
          end 
          if(_th_myfunc_start[12] && (th_blink == 10)) begin
            _th_myfunc_12_tid_309 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[12]) begin
            th_myfunc_12 <= th_myfunc_12_1;
          end 
        end
        th_myfunc_12_1: begin
          _th_myfunc_12_tid_310 <= _th_myfunc_12_tid_309;
          th_myfunc_12 <= th_myfunc_12_2;
        end
        th_myfunc_12_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 12)) begin
            th_myfunc_12 <= th_myfunc_12_3;
          end 
        end
        th_myfunc_12_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 12))) begin
            th_myfunc_12 <= th_myfunc_12_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 12)) begin
            th_myfunc_12 <= th_myfunc_12_4;
          end 
        end
        th_myfunc_12_4: begin
          $display("Thread %d Lock", _th_myfunc_12_tid_310);
          th_myfunc_12 <= th_myfunc_12_5;
        end
        th_myfunc_12_5: begin
          _th_myfunc_12_time_311 <= sw;
          th_myfunc_12 <= th_myfunc_12_6;
        end
        th_myfunc_12_6: begin
          _th_myfunc_12_i_312 <= 0;
          th_myfunc_12 <= th_myfunc_12_7;
        end
        th_myfunc_12_7: begin
          if(_th_myfunc_12_i_312 < _th_myfunc_12_time_311) begin
            th_myfunc_12 <= th_myfunc_12_8;
          end else begin
            th_myfunc_12 <= th_myfunc_12_9;
          end
        end
        th_myfunc_12_8: begin
          _th_myfunc_12_i_312 <= _th_myfunc_12_i_312 + 1;
          th_myfunc_12 <= th_myfunc_12_7;
        end
        th_myfunc_12_9: begin
          th_myfunc_12 <= th_myfunc_12_10;
        end
        th_myfunc_12_10: begin
          $display("Thread %d count = %d", _th_myfunc_12_tid_310, count);
          th_myfunc_12 <= th_myfunc_12_11;
        end
        th_myfunc_12_11: begin
          th_myfunc_12 <= th_myfunc_12_12;
        end
        th_myfunc_12_12: begin
          $display("Thread %d Unlock", _th_myfunc_12_tid_310);
          th_myfunc_12 <= th_myfunc_12_13;
        end
        th_myfunc_12_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 12)) begin
            _th_myfunc_12_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 12)) begin
            th_myfunc_12 <= th_myfunc_12_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_13_1 = 1;
  localparam th_myfunc_13_2 = 2;
  localparam th_myfunc_13_3 = 3;
  localparam th_myfunc_13_4 = 4;
  localparam th_myfunc_13_5 = 5;
  localparam th_myfunc_13_6 = 6;
  localparam th_myfunc_13_7 = 7;
  localparam th_myfunc_13_8 = 8;
  localparam th_myfunc_13_9 = 9;
  localparam th_myfunc_13_10 = 10;
  localparam th_myfunc_13_11 = 11;
  localparam th_myfunc_13_12 = 12;
  localparam th_myfunc_13_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_13 <= th_myfunc_13_init;
      _th_myfunc_13_called <= 0;
      _th_myfunc_13_tid_313 <= 0;
      _th_myfunc_13_tid_314 <= 0;
      _th_myfunc_13_time_315 <= 0;
      _th_myfunc_13_i_316 <= 0;
    end else begin
      case(th_myfunc_13)
        th_myfunc_13_init: begin
          if(_th_myfunc_start[13] && (th_blink == 10)) begin
            _th_myfunc_13_called <= 1;
          end 
          if(_th_myfunc_start[13] && (th_blink == 10)) begin
            _th_myfunc_13_tid_313 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[13]) begin
            th_myfunc_13 <= th_myfunc_13_1;
          end 
        end
        th_myfunc_13_1: begin
          _th_myfunc_13_tid_314 <= _th_myfunc_13_tid_313;
          th_myfunc_13 <= th_myfunc_13_2;
        end
        th_myfunc_13_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 13)) begin
            th_myfunc_13 <= th_myfunc_13_3;
          end 
        end
        th_myfunc_13_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 13))) begin
            th_myfunc_13 <= th_myfunc_13_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 13)) begin
            th_myfunc_13 <= th_myfunc_13_4;
          end 
        end
        th_myfunc_13_4: begin
          $display("Thread %d Lock", _th_myfunc_13_tid_314);
          th_myfunc_13 <= th_myfunc_13_5;
        end
        th_myfunc_13_5: begin
          _th_myfunc_13_time_315 <= sw;
          th_myfunc_13 <= th_myfunc_13_6;
        end
        th_myfunc_13_6: begin
          _th_myfunc_13_i_316 <= 0;
          th_myfunc_13 <= th_myfunc_13_7;
        end
        th_myfunc_13_7: begin
          if(_th_myfunc_13_i_316 < _th_myfunc_13_time_315) begin
            th_myfunc_13 <= th_myfunc_13_8;
          end else begin
            th_myfunc_13 <= th_myfunc_13_9;
          end
        end
        th_myfunc_13_8: begin
          _th_myfunc_13_i_316 <= _th_myfunc_13_i_316 + 1;
          th_myfunc_13 <= th_myfunc_13_7;
        end
        th_myfunc_13_9: begin
          th_myfunc_13 <= th_myfunc_13_10;
        end
        th_myfunc_13_10: begin
          $display("Thread %d count = %d", _th_myfunc_13_tid_314, count);
          th_myfunc_13 <= th_myfunc_13_11;
        end
        th_myfunc_13_11: begin
          th_myfunc_13 <= th_myfunc_13_12;
        end
        th_myfunc_13_12: begin
          $display("Thread %d Unlock", _th_myfunc_13_tid_314);
          th_myfunc_13 <= th_myfunc_13_13;
        end
        th_myfunc_13_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 13)) begin
            _th_myfunc_13_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 13)) begin
            th_myfunc_13 <= th_myfunc_13_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_14_1 = 1;
  localparam th_myfunc_14_2 = 2;
  localparam th_myfunc_14_3 = 3;
  localparam th_myfunc_14_4 = 4;
  localparam th_myfunc_14_5 = 5;
  localparam th_myfunc_14_6 = 6;
  localparam th_myfunc_14_7 = 7;
  localparam th_myfunc_14_8 = 8;
  localparam th_myfunc_14_9 = 9;
  localparam th_myfunc_14_10 = 10;
  localparam th_myfunc_14_11 = 11;
  localparam th_myfunc_14_12 = 12;
  localparam th_myfunc_14_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_14 <= th_myfunc_14_init;
      _th_myfunc_14_called <= 0;
      _th_myfunc_14_tid_317 <= 0;
      _th_myfunc_14_tid_318 <= 0;
      _th_myfunc_14_time_319 <= 0;
      _th_myfunc_14_i_320 <= 0;
    end else begin
      case(th_myfunc_14)
        th_myfunc_14_init: begin
          if(_th_myfunc_start[14] && (th_blink == 10)) begin
            _th_myfunc_14_called <= 1;
          end 
          if(_th_myfunc_start[14] && (th_blink == 10)) begin
            _th_myfunc_14_tid_317 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[14]) begin
            th_myfunc_14 <= th_myfunc_14_1;
          end 
        end
        th_myfunc_14_1: begin
          _th_myfunc_14_tid_318 <= _th_myfunc_14_tid_317;
          th_myfunc_14 <= th_myfunc_14_2;
        end
        th_myfunc_14_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 14)) begin
            th_myfunc_14 <= th_myfunc_14_3;
          end 
        end
        th_myfunc_14_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 14))) begin
            th_myfunc_14 <= th_myfunc_14_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 14)) begin
            th_myfunc_14 <= th_myfunc_14_4;
          end 
        end
        th_myfunc_14_4: begin
          $display("Thread %d Lock", _th_myfunc_14_tid_318);
          th_myfunc_14 <= th_myfunc_14_5;
        end
        th_myfunc_14_5: begin
          _th_myfunc_14_time_319 <= sw;
          th_myfunc_14 <= th_myfunc_14_6;
        end
        th_myfunc_14_6: begin
          _th_myfunc_14_i_320 <= 0;
          th_myfunc_14 <= th_myfunc_14_7;
        end
        th_myfunc_14_7: begin
          if(_th_myfunc_14_i_320 < _th_myfunc_14_time_319) begin
            th_myfunc_14 <= th_myfunc_14_8;
          end else begin
            th_myfunc_14 <= th_myfunc_14_9;
          end
        end
        th_myfunc_14_8: begin
          _th_myfunc_14_i_320 <= _th_myfunc_14_i_320 + 1;
          th_myfunc_14 <= th_myfunc_14_7;
        end
        th_myfunc_14_9: begin
          th_myfunc_14 <= th_myfunc_14_10;
        end
        th_myfunc_14_10: begin
          $display("Thread %d count = %d", _th_myfunc_14_tid_318, count);
          th_myfunc_14 <= th_myfunc_14_11;
        end
        th_myfunc_14_11: begin
          th_myfunc_14 <= th_myfunc_14_12;
        end
        th_myfunc_14_12: begin
          $display("Thread %d Unlock", _th_myfunc_14_tid_318);
          th_myfunc_14 <= th_myfunc_14_13;
        end
        th_myfunc_14_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 14)) begin
            _th_myfunc_14_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 14)) begin
            th_myfunc_14 <= th_myfunc_14_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_15_1 = 1;
  localparam th_myfunc_15_2 = 2;
  localparam th_myfunc_15_3 = 3;
  localparam th_myfunc_15_4 = 4;
  localparam th_myfunc_15_5 = 5;
  localparam th_myfunc_15_6 = 6;
  localparam th_myfunc_15_7 = 7;
  localparam th_myfunc_15_8 = 8;
  localparam th_myfunc_15_9 = 9;
  localparam th_myfunc_15_10 = 10;
  localparam th_myfunc_15_11 = 11;
  localparam th_myfunc_15_12 = 12;
  localparam th_myfunc_15_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_15 <= th_myfunc_15_init;
      _th_myfunc_15_called <= 0;
      _th_myfunc_15_tid_321 <= 0;
      _th_myfunc_15_tid_322 <= 0;
      _th_myfunc_15_time_323 <= 0;
      _th_myfunc_15_i_324 <= 0;
    end else begin
      case(th_myfunc_15)
        th_myfunc_15_init: begin
          if(_th_myfunc_start[15] && (th_blink == 10)) begin
            _th_myfunc_15_called <= 1;
          end 
          if(_th_myfunc_start[15] && (th_blink == 10)) begin
            _th_myfunc_15_tid_321 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[15]) begin
            th_myfunc_15 <= th_myfunc_15_1;
          end 
        end
        th_myfunc_15_1: begin
          _th_myfunc_15_tid_322 <= _th_myfunc_15_tid_321;
          th_myfunc_15 <= th_myfunc_15_2;
        end
        th_myfunc_15_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 15)) begin
            th_myfunc_15 <= th_myfunc_15_3;
          end 
        end
        th_myfunc_15_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 15))) begin
            th_myfunc_15 <= th_myfunc_15_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 15)) begin
            th_myfunc_15 <= th_myfunc_15_4;
          end 
        end
        th_myfunc_15_4: begin
          $display("Thread %d Lock", _th_myfunc_15_tid_322);
          th_myfunc_15 <= th_myfunc_15_5;
        end
        th_myfunc_15_5: begin
          _th_myfunc_15_time_323 <= sw;
          th_myfunc_15 <= th_myfunc_15_6;
        end
        th_myfunc_15_6: begin
          _th_myfunc_15_i_324 <= 0;
          th_myfunc_15 <= th_myfunc_15_7;
        end
        th_myfunc_15_7: begin
          if(_th_myfunc_15_i_324 < _th_myfunc_15_time_323) begin
            th_myfunc_15 <= th_myfunc_15_8;
          end else begin
            th_myfunc_15 <= th_myfunc_15_9;
          end
        end
        th_myfunc_15_8: begin
          _th_myfunc_15_i_324 <= _th_myfunc_15_i_324 + 1;
          th_myfunc_15 <= th_myfunc_15_7;
        end
        th_myfunc_15_9: begin
          th_myfunc_15 <= th_myfunc_15_10;
        end
        th_myfunc_15_10: begin
          $display("Thread %d count = %d", _th_myfunc_15_tid_322, count);
          th_myfunc_15 <= th_myfunc_15_11;
        end
        th_myfunc_15_11: begin
          th_myfunc_15 <= th_myfunc_15_12;
        end
        th_myfunc_15_12: begin
          $display("Thread %d Unlock", _th_myfunc_15_tid_322);
          th_myfunc_15 <= th_myfunc_15_13;
        end
        th_myfunc_15_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 15)) begin
            _th_myfunc_15_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 15)) begin
            th_myfunc_15 <= th_myfunc_15_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_16_1 = 1;
  localparam th_myfunc_16_2 = 2;
  localparam th_myfunc_16_3 = 3;
  localparam th_myfunc_16_4 = 4;
  localparam th_myfunc_16_5 = 5;
  localparam th_myfunc_16_6 = 6;
  localparam th_myfunc_16_7 = 7;
  localparam th_myfunc_16_8 = 8;
  localparam th_myfunc_16_9 = 9;
  localparam th_myfunc_16_10 = 10;
  localparam th_myfunc_16_11 = 11;
  localparam th_myfunc_16_12 = 12;
  localparam th_myfunc_16_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_16 <= th_myfunc_16_init;
      _th_myfunc_16_called <= 0;
      _th_myfunc_16_tid_325 <= 0;
      _th_myfunc_16_tid_326 <= 0;
      _th_myfunc_16_time_327 <= 0;
      _th_myfunc_16_i_328 <= 0;
    end else begin
      case(th_myfunc_16)
        th_myfunc_16_init: begin
          if(_th_myfunc_start[16] && (th_blink == 10)) begin
            _th_myfunc_16_called <= 1;
          end 
          if(_th_myfunc_start[16] && (th_blink == 10)) begin
            _th_myfunc_16_tid_325 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[16]) begin
            th_myfunc_16 <= th_myfunc_16_1;
          end 
        end
        th_myfunc_16_1: begin
          _th_myfunc_16_tid_326 <= _th_myfunc_16_tid_325;
          th_myfunc_16 <= th_myfunc_16_2;
        end
        th_myfunc_16_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 16)) begin
            th_myfunc_16 <= th_myfunc_16_3;
          end 
        end
        th_myfunc_16_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 16))) begin
            th_myfunc_16 <= th_myfunc_16_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 16)) begin
            th_myfunc_16 <= th_myfunc_16_4;
          end 
        end
        th_myfunc_16_4: begin
          $display("Thread %d Lock", _th_myfunc_16_tid_326);
          th_myfunc_16 <= th_myfunc_16_5;
        end
        th_myfunc_16_5: begin
          _th_myfunc_16_time_327 <= sw;
          th_myfunc_16 <= th_myfunc_16_6;
        end
        th_myfunc_16_6: begin
          _th_myfunc_16_i_328 <= 0;
          th_myfunc_16 <= th_myfunc_16_7;
        end
        th_myfunc_16_7: begin
          if(_th_myfunc_16_i_328 < _th_myfunc_16_time_327) begin
            th_myfunc_16 <= th_myfunc_16_8;
          end else begin
            th_myfunc_16 <= th_myfunc_16_9;
          end
        end
        th_myfunc_16_8: begin
          _th_myfunc_16_i_328 <= _th_myfunc_16_i_328 + 1;
          th_myfunc_16 <= th_myfunc_16_7;
        end
        th_myfunc_16_9: begin
          th_myfunc_16 <= th_myfunc_16_10;
        end
        th_myfunc_16_10: begin
          $display("Thread %d count = %d", _th_myfunc_16_tid_326, count);
          th_myfunc_16 <= th_myfunc_16_11;
        end
        th_myfunc_16_11: begin
          th_myfunc_16 <= th_myfunc_16_12;
        end
        th_myfunc_16_12: begin
          $display("Thread %d Unlock", _th_myfunc_16_tid_326);
          th_myfunc_16 <= th_myfunc_16_13;
        end
        th_myfunc_16_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 16)) begin
            _th_myfunc_16_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 16)) begin
            th_myfunc_16 <= th_myfunc_16_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_17_1 = 1;
  localparam th_myfunc_17_2 = 2;
  localparam th_myfunc_17_3 = 3;
  localparam th_myfunc_17_4 = 4;
  localparam th_myfunc_17_5 = 5;
  localparam th_myfunc_17_6 = 6;
  localparam th_myfunc_17_7 = 7;
  localparam th_myfunc_17_8 = 8;
  localparam th_myfunc_17_9 = 9;
  localparam th_myfunc_17_10 = 10;
  localparam th_myfunc_17_11 = 11;
  localparam th_myfunc_17_12 = 12;
  localparam th_myfunc_17_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_17 <= th_myfunc_17_init;
      _th_myfunc_17_called <= 0;
      _th_myfunc_17_tid_329 <= 0;
      _th_myfunc_17_tid_330 <= 0;
      _th_myfunc_17_time_331 <= 0;
      _th_myfunc_17_i_332 <= 0;
    end else begin
      case(th_myfunc_17)
        th_myfunc_17_init: begin
          if(_th_myfunc_start[17] && (th_blink == 10)) begin
            _th_myfunc_17_called <= 1;
          end 
          if(_th_myfunc_start[17] && (th_blink == 10)) begin
            _th_myfunc_17_tid_329 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[17]) begin
            th_myfunc_17 <= th_myfunc_17_1;
          end 
        end
        th_myfunc_17_1: begin
          _th_myfunc_17_tid_330 <= _th_myfunc_17_tid_329;
          th_myfunc_17 <= th_myfunc_17_2;
        end
        th_myfunc_17_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 17)) begin
            th_myfunc_17 <= th_myfunc_17_3;
          end 
        end
        th_myfunc_17_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 17))) begin
            th_myfunc_17 <= th_myfunc_17_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 17)) begin
            th_myfunc_17 <= th_myfunc_17_4;
          end 
        end
        th_myfunc_17_4: begin
          $display("Thread %d Lock", _th_myfunc_17_tid_330);
          th_myfunc_17 <= th_myfunc_17_5;
        end
        th_myfunc_17_5: begin
          _th_myfunc_17_time_331 <= sw;
          th_myfunc_17 <= th_myfunc_17_6;
        end
        th_myfunc_17_6: begin
          _th_myfunc_17_i_332 <= 0;
          th_myfunc_17 <= th_myfunc_17_7;
        end
        th_myfunc_17_7: begin
          if(_th_myfunc_17_i_332 < _th_myfunc_17_time_331) begin
            th_myfunc_17 <= th_myfunc_17_8;
          end else begin
            th_myfunc_17 <= th_myfunc_17_9;
          end
        end
        th_myfunc_17_8: begin
          _th_myfunc_17_i_332 <= _th_myfunc_17_i_332 + 1;
          th_myfunc_17 <= th_myfunc_17_7;
        end
        th_myfunc_17_9: begin
          th_myfunc_17 <= th_myfunc_17_10;
        end
        th_myfunc_17_10: begin
          $display("Thread %d count = %d", _th_myfunc_17_tid_330, count);
          th_myfunc_17 <= th_myfunc_17_11;
        end
        th_myfunc_17_11: begin
          th_myfunc_17 <= th_myfunc_17_12;
        end
        th_myfunc_17_12: begin
          $display("Thread %d Unlock", _th_myfunc_17_tid_330);
          th_myfunc_17 <= th_myfunc_17_13;
        end
        th_myfunc_17_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 17)) begin
            _th_myfunc_17_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 17)) begin
            th_myfunc_17 <= th_myfunc_17_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_18_1 = 1;
  localparam th_myfunc_18_2 = 2;
  localparam th_myfunc_18_3 = 3;
  localparam th_myfunc_18_4 = 4;
  localparam th_myfunc_18_5 = 5;
  localparam th_myfunc_18_6 = 6;
  localparam th_myfunc_18_7 = 7;
  localparam th_myfunc_18_8 = 8;
  localparam th_myfunc_18_9 = 9;
  localparam th_myfunc_18_10 = 10;
  localparam th_myfunc_18_11 = 11;
  localparam th_myfunc_18_12 = 12;
  localparam th_myfunc_18_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_18 <= th_myfunc_18_init;
      _th_myfunc_18_called <= 0;
      _th_myfunc_18_tid_333 <= 0;
      _th_myfunc_18_tid_334 <= 0;
      _th_myfunc_18_time_335 <= 0;
      _th_myfunc_18_i_336 <= 0;
    end else begin
      case(th_myfunc_18)
        th_myfunc_18_init: begin
          if(_th_myfunc_start[18] && (th_blink == 10)) begin
            _th_myfunc_18_called <= 1;
          end 
          if(_th_myfunc_start[18] && (th_blink == 10)) begin
            _th_myfunc_18_tid_333 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[18]) begin
            th_myfunc_18 <= th_myfunc_18_1;
          end 
        end
        th_myfunc_18_1: begin
          _th_myfunc_18_tid_334 <= _th_myfunc_18_tid_333;
          th_myfunc_18 <= th_myfunc_18_2;
        end
        th_myfunc_18_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 18)) begin
            th_myfunc_18 <= th_myfunc_18_3;
          end 
        end
        th_myfunc_18_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 18))) begin
            th_myfunc_18 <= th_myfunc_18_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 18)) begin
            th_myfunc_18 <= th_myfunc_18_4;
          end 
        end
        th_myfunc_18_4: begin
          $display("Thread %d Lock", _th_myfunc_18_tid_334);
          th_myfunc_18 <= th_myfunc_18_5;
        end
        th_myfunc_18_5: begin
          _th_myfunc_18_time_335 <= sw;
          th_myfunc_18 <= th_myfunc_18_6;
        end
        th_myfunc_18_6: begin
          _th_myfunc_18_i_336 <= 0;
          th_myfunc_18 <= th_myfunc_18_7;
        end
        th_myfunc_18_7: begin
          if(_th_myfunc_18_i_336 < _th_myfunc_18_time_335) begin
            th_myfunc_18 <= th_myfunc_18_8;
          end else begin
            th_myfunc_18 <= th_myfunc_18_9;
          end
        end
        th_myfunc_18_8: begin
          _th_myfunc_18_i_336 <= _th_myfunc_18_i_336 + 1;
          th_myfunc_18 <= th_myfunc_18_7;
        end
        th_myfunc_18_9: begin
          th_myfunc_18 <= th_myfunc_18_10;
        end
        th_myfunc_18_10: begin
          $display("Thread %d count = %d", _th_myfunc_18_tid_334, count);
          th_myfunc_18 <= th_myfunc_18_11;
        end
        th_myfunc_18_11: begin
          th_myfunc_18 <= th_myfunc_18_12;
        end
        th_myfunc_18_12: begin
          $display("Thread %d Unlock", _th_myfunc_18_tid_334);
          th_myfunc_18 <= th_myfunc_18_13;
        end
        th_myfunc_18_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 18)) begin
            _th_myfunc_18_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 18)) begin
            th_myfunc_18 <= th_myfunc_18_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_19_1 = 1;
  localparam th_myfunc_19_2 = 2;
  localparam th_myfunc_19_3 = 3;
  localparam th_myfunc_19_4 = 4;
  localparam th_myfunc_19_5 = 5;
  localparam th_myfunc_19_6 = 6;
  localparam th_myfunc_19_7 = 7;
  localparam th_myfunc_19_8 = 8;
  localparam th_myfunc_19_9 = 9;
  localparam th_myfunc_19_10 = 10;
  localparam th_myfunc_19_11 = 11;
  localparam th_myfunc_19_12 = 12;
  localparam th_myfunc_19_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_19 <= th_myfunc_19_init;
      _th_myfunc_19_called <= 0;
      _th_myfunc_19_tid_337 <= 0;
      _th_myfunc_19_tid_338 <= 0;
      _th_myfunc_19_time_339 <= 0;
      _th_myfunc_19_i_340 <= 0;
    end else begin
      case(th_myfunc_19)
        th_myfunc_19_init: begin
          if(_th_myfunc_start[19] && (th_blink == 10)) begin
            _th_myfunc_19_called <= 1;
          end 
          if(_th_myfunc_start[19] && (th_blink == 10)) begin
            _th_myfunc_19_tid_337 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[19]) begin
            th_myfunc_19 <= th_myfunc_19_1;
          end 
        end
        th_myfunc_19_1: begin
          _th_myfunc_19_tid_338 <= _th_myfunc_19_tid_337;
          th_myfunc_19 <= th_myfunc_19_2;
        end
        th_myfunc_19_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 19)) begin
            th_myfunc_19 <= th_myfunc_19_3;
          end 
        end
        th_myfunc_19_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 19))) begin
            th_myfunc_19 <= th_myfunc_19_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 19)) begin
            th_myfunc_19 <= th_myfunc_19_4;
          end 
        end
        th_myfunc_19_4: begin
          $display("Thread %d Lock", _th_myfunc_19_tid_338);
          th_myfunc_19 <= th_myfunc_19_5;
        end
        th_myfunc_19_5: begin
          _th_myfunc_19_time_339 <= sw;
          th_myfunc_19 <= th_myfunc_19_6;
        end
        th_myfunc_19_6: begin
          _th_myfunc_19_i_340 <= 0;
          th_myfunc_19 <= th_myfunc_19_7;
        end
        th_myfunc_19_7: begin
          if(_th_myfunc_19_i_340 < _th_myfunc_19_time_339) begin
            th_myfunc_19 <= th_myfunc_19_8;
          end else begin
            th_myfunc_19 <= th_myfunc_19_9;
          end
        end
        th_myfunc_19_8: begin
          _th_myfunc_19_i_340 <= _th_myfunc_19_i_340 + 1;
          th_myfunc_19 <= th_myfunc_19_7;
        end
        th_myfunc_19_9: begin
          th_myfunc_19 <= th_myfunc_19_10;
        end
        th_myfunc_19_10: begin
          $display("Thread %d count = %d", _th_myfunc_19_tid_338, count);
          th_myfunc_19 <= th_myfunc_19_11;
        end
        th_myfunc_19_11: begin
          th_myfunc_19 <= th_myfunc_19_12;
        end
        th_myfunc_19_12: begin
          $display("Thread %d Unlock", _th_myfunc_19_tid_338);
          th_myfunc_19 <= th_myfunc_19_13;
        end
        th_myfunc_19_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 19)) begin
            _th_myfunc_19_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 19)) begin
            th_myfunc_19 <= th_myfunc_19_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_20_1 = 1;
  localparam th_myfunc_20_2 = 2;
  localparam th_myfunc_20_3 = 3;
  localparam th_myfunc_20_4 = 4;
  localparam th_myfunc_20_5 = 5;
  localparam th_myfunc_20_6 = 6;
  localparam th_myfunc_20_7 = 7;
  localparam th_myfunc_20_8 = 8;
  localparam th_myfunc_20_9 = 9;
  localparam th_myfunc_20_10 = 10;
  localparam th_myfunc_20_11 = 11;
  localparam th_myfunc_20_12 = 12;
  localparam th_myfunc_20_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_20 <= th_myfunc_20_init;
      _th_myfunc_20_called <= 0;
      _th_myfunc_20_tid_341 <= 0;
      _th_myfunc_20_tid_342 <= 0;
      _th_myfunc_20_time_343 <= 0;
      _th_myfunc_20_i_344 <= 0;
    end else begin
      case(th_myfunc_20)
        th_myfunc_20_init: begin
          if(_th_myfunc_start[20] && (th_blink == 10)) begin
            _th_myfunc_20_called <= 1;
          end 
          if(_th_myfunc_start[20] && (th_blink == 10)) begin
            _th_myfunc_20_tid_341 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[20]) begin
            th_myfunc_20 <= th_myfunc_20_1;
          end 
        end
        th_myfunc_20_1: begin
          _th_myfunc_20_tid_342 <= _th_myfunc_20_tid_341;
          th_myfunc_20 <= th_myfunc_20_2;
        end
        th_myfunc_20_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 20)) begin
            th_myfunc_20 <= th_myfunc_20_3;
          end 
        end
        th_myfunc_20_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 20))) begin
            th_myfunc_20 <= th_myfunc_20_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 20)) begin
            th_myfunc_20 <= th_myfunc_20_4;
          end 
        end
        th_myfunc_20_4: begin
          $display("Thread %d Lock", _th_myfunc_20_tid_342);
          th_myfunc_20 <= th_myfunc_20_5;
        end
        th_myfunc_20_5: begin
          _th_myfunc_20_time_343 <= sw;
          th_myfunc_20 <= th_myfunc_20_6;
        end
        th_myfunc_20_6: begin
          _th_myfunc_20_i_344 <= 0;
          th_myfunc_20 <= th_myfunc_20_7;
        end
        th_myfunc_20_7: begin
          if(_th_myfunc_20_i_344 < _th_myfunc_20_time_343) begin
            th_myfunc_20 <= th_myfunc_20_8;
          end else begin
            th_myfunc_20 <= th_myfunc_20_9;
          end
        end
        th_myfunc_20_8: begin
          _th_myfunc_20_i_344 <= _th_myfunc_20_i_344 + 1;
          th_myfunc_20 <= th_myfunc_20_7;
        end
        th_myfunc_20_9: begin
          th_myfunc_20 <= th_myfunc_20_10;
        end
        th_myfunc_20_10: begin
          $display("Thread %d count = %d", _th_myfunc_20_tid_342, count);
          th_myfunc_20 <= th_myfunc_20_11;
        end
        th_myfunc_20_11: begin
          th_myfunc_20 <= th_myfunc_20_12;
        end
        th_myfunc_20_12: begin
          $display("Thread %d Unlock", _th_myfunc_20_tid_342);
          th_myfunc_20 <= th_myfunc_20_13;
        end
        th_myfunc_20_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 20)) begin
            _th_myfunc_20_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 20)) begin
            th_myfunc_20 <= th_myfunc_20_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_21_1 = 1;
  localparam th_myfunc_21_2 = 2;
  localparam th_myfunc_21_3 = 3;
  localparam th_myfunc_21_4 = 4;
  localparam th_myfunc_21_5 = 5;
  localparam th_myfunc_21_6 = 6;
  localparam th_myfunc_21_7 = 7;
  localparam th_myfunc_21_8 = 8;
  localparam th_myfunc_21_9 = 9;
  localparam th_myfunc_21_10 = 10;
  localparam th_myfunc_21_11 = 11;
  localparam th_myfunc_21_12 = 12;
  localparam th_myfunc_21_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_21 <= th_myfunc_21_init;
      _th_myfunc_21_called <= 0;
      _th_myfunc_21_tid_345 <= 0;
      _th_myfunc_21_tid_346 <= 0;
      _th_myfunc_21_time_347 <= 0;
      _th_myfunc_21_i_348 <= 0;
    end else begin
      case(th_myfunc_21)
        th_myfunc_21_init: begin
          if(_th_myfunc_start[21] && (th_blink == 10)) begin
            _th_myfunc_21_called <= 1;
          end 
          if(_th_myfunc_start[21] && (th_blink == 10)) begin
            _th_myfunc_21_tid_345 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[21]) begin
            th_myfunc_21 <= th_myfunc_21_1;
          end 
        end
        th_myfunc_21_1: begin
          _th_myfunc_21_tid_346 <= _th_myfunc_21_tid_345;
          th_myfunc_21 <= th_myfunc_21_2;
        end
        th_myfunc_21_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 21)) begin
            th_myfunc_21 <= th_myfunc_21_3;
          end 
        end
        th_myfunc_21_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 21))) begin
            th_myfunc_21 <= th_myfunc_21_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 21)) begin
            th_myfunc_21 <= th_myfunc_21_4;
          end 
        end
        th_myfunc_21_4: begin
          $display("Thread %d Lock", _th_myfunc_21_tid_346);
          th_myfunc_21 <= th_myfunc_21_5;
        end
        th_myfunc_21_5: begin
          _th_myfunc_21_time_347 <= sw;
          th_myfunc_21 <= th_myfunc_21_6;
        end
        th_myfunc_21_6: begin
          _th_myfunc_21_i_348 <= 0;
          th_myfunc_21 <= th_myfunc_21_7;
        end
        th_myfunc_21_7: begin
          if(_th_myfunc_21_i_348 < _th_myfunc_21_time_347) begin
            th_myfunc_21 <= th_myfunc_21_8;
          end else begin
            th_myfunc_21 <= th_myfunc_21_9;
          end
        end
        th_myfunc_21_8: begin
          _th_myfunc_21_i_348 <= _th_myfunc_21_i_348 + 1;
          th_myfunc_21 <= th_myfunc_21_7;
        end
        th_myfunc_21_9: begin
          th_myfunc_21 <= th_myfunc_21_10;
        end
        th_myfunc_21_10: begin
          $display("Thread %d count = %d", _th_myfunc_21_tid_346, count);
          th_myfunc_21 <= th_myfunc_21_11;
        end
        th_myfunc_21_11: begin
          th_myfunc_21 <= th_myfunc_21_12;
        end
        th_myfunc_21_12: begin
          $display("Thread %d Unlock", _th_myfunc_21_tid_346);
          th_myfunc_21 <= th_myfunc_21_13;
        end
        th_myfunc_21_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 21)) begin
            _th_myfunc_21_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 21)) begin
            th_myfunc_21 <= th_myfunc_21_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_22_1 = 1;
  localparam th_myfunc_22_2 = 2;
  localparam th_myfunc_22_3 = 3;
  localparam th_myfunc_22_4 = 4;
  localparam th_myfunc_22_5 = 5;
  localparam th_myfunc_22_6 = 6;
  localparam th_myfunc_22_7 = 7;
  localparam th_myfunc_22_8 = 8;
  localparam th_myfunc_22_9 = 9;
  localparam th_myfunc_22_10 = 10;
  localparam th_myfunc_22_11 = 11;
  localparam th_myfunc_22_12 = 12;
  localparam th_myfunc_22_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_22 <= th_myfunc_22_init;
      _th_myfunc_22_called <= 0;
      _th_myfunc_22_tid_349 <= 0;
      _th_myfunc_22_tid_350 <= 0;
      _th_myfunc_22_time_351 <= 0;
      _th_myfunc_22_i_352 <= 0;
    end else begin
      case(th_myfunc_22)
        th_myfunc_22_init: begin
          if(_th_myfunc_start[22] && (th_blink == 10)) begin
            _th_myfunc_22_called <= 1;
          end 
          if(_th_myfunc_start[22] && (th_blink == 10)) begin
            _th_myfunc_22_tid_349 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[22]) begin
            th_myfunc_22 <= th_myfunc_22_1;
          end 
        end
        th_myfunc_22_1: begin
          _th_myfunc_22_tid_350 <= _th_myfunc_22_tid_349;
          th_myfunc_22 <= th_myfunc_22_2;
        end
        th_myfunc_22_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 22)) begin
            th_myfunc_22 <= th_myfunc_22_3;
          end 
        end
        th_myfunc_22_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 22))) begin
            th_myfunc_22 <= th_myfunc_22_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 22)) begin
            th_myfunc_22 <= th_myfunc_22_4;
          end 
        end
        th_myfunc_22_4: begin
          $display("Thread %d Lock", _th_myfunc_22_tid_350);
          th_myfunc_22 <= th_myfunc_22_5;
        end
        th_myfunc_22_5: begin
          _th_myfunc_22_time_351 <= sw;
          th_myfunc_22 <= th_myfunc_22_6;
        end
        th_myfunc_22_6: begin
          _th_myfunc_22_i_352 <= 0;
          th_myfunc_22 <= th_myfunc_22_7;
        end
        th_myfunc_22_7: begin
          if(_th_myfunc_22_i_352 < _th_myfunc_22_time_351) begin
            th_myfunc_22 <= th_myfunc_22_8;
          end else begin
            th_myfunc_22 <= th_myfunc_22_9;
          end
        end
        th_myfunc_22_8: begin
          _th_myfunc_22_i_352 <= _th_myfunc_22_i_352 + 1;
          th_myfunc_22 <= th_myfunc_22_7;
        end
        th_myfunc_22_9: begin
          th_myfunc_22 <= th_myfunc_22_10;
        end
        th_myfunc_22_10: begin
          $display("Thread %d count = %d", _th_myfunc_22_tid_350, count);
          th_myfunc_22 <= th_myfunc_22_11;
        end
        th_myfunc_22_11: begin
          th_myfunc_22 <= th_myfunc_22_12;
        end
        th_myfunc_22_12: begin
          $display("Thread %d Unlock", _th_myfunc_22_tid_350);
          th_myfunc_22 <= th_myfunc_22_13;
        end
        th_myfunc_22_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 22)) begin
            _th_myfunc_22_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 22)) begin
            th_myfunc_22 <= th_myfunc_22_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_23_1 = 1;
  localparam th_myfunc_23_2 = 2;
  localparam th_myfunc_23_3 = 3;
  localparam th_myfunc_23_4 = 4;
  localparam th_myfunc_23_5 = 5;
  localparam th_myfunc_23_6 = 6;
  localparam th_myfunc_23_7 = 7;
  localparam th_myfunc_23_8 = 8;
  localparam th_myfunc_23_9 = 9;
  localparam th_myfunc_23_10 = 10;
  localparam th_myfunc_23_11 = 11;
  localparam th_myfunc_23_12 = 12;
  localparam th_myfunc_23_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_23 <= th_myfunc_23_init;
      _th_myfunc_23_called <= 0;
      _th_myfunc_23_tid_353 <= 0;
      _th_myfunc_23_tid_354 <= 0;
      _th_myfunc_23_time_355 <= 0;
      _th_myfunc_23_i_356 <= 0;
    end else begin
      case(th_myfunc_23)
        th_myfunc_23_init: begin
          if(_th_myfunc_start[23] && (th_blink == 10)) begin
            _th_myfunc_23_called <= 1;
          end 
          if(_th_myfunc_start[23] && (th_blink == 10)) begin
            _th_myfunc_23_tid_353 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[23]) begin
            th_myfunc_23 <= th_myfunc_23_1;
          end 
        end
        th_myfunc_23_1: begin
          _th_myfunc_23_tid_354 <= _th_myfunc_23_tid_353;
          th_myfunc_23 <= th_myfunc_23_2;
        end
        th_myfunc_23_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 23)) begin
            th_myfunc_23 <= th_myfunc_23_3;
          end 
        end
        th_myfunc_23_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 23))) begin
            th_myfunc_23 <= th_myfunc_23_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 23)) begin
            th_myfunc_23 <= th_myfunc_23_4;
          end 
        end
        th_myfunc_23_4: begin
          $display("Thread %d Lock", _th_myfunc_23_tid_354);
          th_myfunc_23 <= th_myfunc_23_5;
        end
        th_myfunc_23_5: begin
          _th_myfunc_23_time_355 <= sw;
          th_myfunc_23 <= th_myfunc_23_6;
        end
        th_myfunc_23_6: begin
          _th_myfunc_23_i_356 <= 0;
          th_myfunc_23 <= th_myfunc_23_7;
        end
        th_myfunc_23_7: begin
          if(_th_myfunc_23_i_356 < _th_myfunc_23_time_355) begin
            th_myfunc_23 <= th_myfunc_23_8;
          end else begin
            th_myfunc_23 <= th_myfunc_23_9;
          end
        end
        th_myfunc_23_8: begin
          _th_myfunc_23_i_356 <= _th_myfunc_23_i_356 + 1;
          th_myfunc_23 <= th_myfunc_23_7;
        end
        th_myfunc_23_9: begin
          th_myfunc_23 <= th_myfunc_23_10;
        end
        th_myfunc_23_10: begin
          $display("Thread %d count = %d", _th_myfunc_23_tid_354, count);
          th_myfunc_23 <= th_myfunc_23_11;
        end
        th_myfunc_23_11: begin
          th_myfunc_23 <= th_myfunc_23_12;
        end
        th_myfunc_23_12: begin
          $display("Thread %d Unlock", _th_myfunc_23_tid_354);
          th_myfunc_23 <= th_myfunc_23_13;
        end
        th_myfunc_23_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 23)) begin
            _th_myfunc_23_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 23)) begin
            th_myfunc_23 <= th_myfunc_23_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_24_1 = 1;
  localparam th_myfunc_24_2 = 2;
  localparam th_myfunc_24_3 = 3;
  localparam th_myfunc_24_4 = 4;
  localparam th_myfunc_24_5 = 5;
  localparam th_myfunc_24_6 = 6;
  localparam th_myfunc_24_7 = 7;
  localparam th_myfunc_24_8 = 8;
  localparam th_myfunc_24_9 = 9;
  localparam th_myfunc_24_10 = 10;
  localparam th_myfunc_24_11 = 11;
  localparam th_myfunc_24_12 = 12;
  localparam th_myfunc_24_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_24 <= th_myfunc_24_init;
      _th_myfunc_24_called <= 0;
      _th_myfunc_24_tid_357 <= 0;
      _th_myfunc_24_tid_358 <= 0;
      _th_myfunc_24_time_359 <= 0;
      _th_myfunc_24_i_360 <= 0;
    end else begin
      case(th_myfunc_24)
        th_myfunc_24_init: begin
          if(_th_myfunc_start[24] && (th_blink == 10)) begin
            _th_myfunc_24_called <= 1;
          end 
          if(_th_myfunc_start[24] && (th_blink == 10)) begin
            _th_myfunc_24_tid_357 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[24]) begin
            th_myfunc_24 <= th_myfunc_24_1;
          end 
        end
        th_myfunc_24_1: begin
          _th_myfunc_24_tid_358 <= _th_myfunc_24_tid_357;
          th_myfunc_24 <= th_myfunc_24_2;
        end
        th_myfunc_24_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 24)) begin
            th_myfunc_24 <= th_myfunc_24_3;
          end 
        end
        th_myfunc_24_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 24))) begin
            th_myfunc_24 <= th_myfunc_24_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 24)) begin
            th_myfunc_24 <= th_myfunc_24_4;
          end 
        end
        th_myfunc_24_4: begin
          $display("Thread %d Lock", _th_myfunc_24_tid_358);
          th_myfunc_24 <= th_myfunc_24_5;
        end
        th_myfunc_24_5: begin
          _th_myfunc_24_time_359 <= sw;
          th_myfunc_24 <= th_myfunc_24_6;
        end
        th_myfunc_24_6: begin
          _th_myfunc_24_i_360 <= 0;
          th_myfunc_24 <= th_myfunc_24_7;
        end
        th_myfunc_24_7: begin
          if(_th_myfunc_24_i_360 < _th_myfunc_24_time_359) begin
            th_myfunc_24 <= th_myfunc_24_8;
          end else begin
            th_myfunc_24 <= th_myfunc_24_9;
          end
        end
        th_myfunc_24_8: begin
          _th_myfunc_24_i_360 <= _th_myfunc_24_i_360 + 1;
          th_myfunc_24 <= th_myfunc_24_7;
        end
        th_myfunc_24_9: begin
          th_myfunc_24 <= th_myfunc_24_10;
        end
        th_myfunc_24_10: begin
          $display("Thread %d count = %d", _th_myfunc_24_tid_358, count);
          th_myfunc_24 <= th_myfunc_24_11;
        end
        th_myfunc_24_11: begin
          th_myfunc_24 <= th_myfunc_24_12;
        end
        th_myfunc_24_12: begin
          $display("Thread %d Unlock", _th_myfunc_24_tid_358);
          th_myfunc_24 <= th_myfunc_24_13;
        end
        th_myfunc_24_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 24)) begin
            _th_myfunc_24_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 24)) begin
            th_myfunc_24 <= th_myfunc_24_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_25_1 = 1;
  localparam th_myfunc_25_2 = 2;
  localparam th_myfunc_25_3 = 3;
  localparam th_myfunc_25_4 = 4;
  localparam th_myfunc_25_5 = 5;
  localparam th_myfunc_25_6 = 6;
  localparam th_myfunc_25_7 = 7;
  localparam th_myfunc_25_8 = 8;
  localparam th_myfunc_25_9 = 9;
  localparam th_myfunc_25_10 = 10;
  localparam th_myfunc_25_11 = 11;
  localparam th_myfunc_25_12 = 12;
  localparam th_myfunc_25_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_25 <= th_myfunc_25_init;
      _th_myfunc_25_called <= 0;
      _th_myfunc_25_tid_361 <= 0;
      _th_myfunc_25_tid_362 <= 0;
      _th_myfunc_25_time_363 <= 0;
      _th_myfunc_25_i_364 <= 0;
    end else begin
      case(th_myfunc_25)
        th_myfunc_25_init: begin
          if(_th_myfunc_start[25] && (th_blink == 10)) begin
            _th_myfunc_25_called <= 1;
          end 
          if(_th_myfunc_start[25] && (th_blink == 10)) begin
            _th_myfunc_25_tid_361 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[25]) begin
            th_myfunc_25 <= th_myfunc_25_1;
          end 
        end
        th_myfunc_25_1: begin
          _th_myfunc_25_tid_362 <= _th_myfunc_25_tid_361;
          th_myfunc_25 <= th_myfunc_25_2;
        end
        th_myfunc_25_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 25)) begin
            th_myfunc_25 <= th_myfunc_25_3;
          end 
        end
        th_myfunc_25_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 25))) begin
            th_myfunc_25 <= th_myfunc_25_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 25)) begin
            th_myfunc_25 <= th_myfunc_25_4;
          end 
        end
        th_myfunc_25_4: begin
          $display("Thread %d Lock", _th_myfunc_25_tid_362);
          th_myfunc_25 <= th_myfunc_25_5;
        end
        th_myfunc_25_5: begin
          _th_myfunc_25_time_363 <= sw;
          th_myfunc_25 <= th_myfunc_25_6;
        end
        th_myfunc_25_6: begin
          _th_myfunc_25_i_364 <= 0;
          th_myfunc_25 <= th_myfunc_25_7;
        end
        th_myfunc_25_7: begin
          if(_th_myfunc_25_i_364 < _th_myfunc_25_time_363) begin
            th_myfunc_25 <= th_myfunc_25_8;
          end else begin
            th_myfunc_25 <= th_myfunc_25_9;
          end
        end
        th_myfunc_25_8: begin
          _th_myfunc_25_i_364 <= _th_myfunc_25_i_364 + 1;
          th_myfunc_25 <= th_myfunc_25_7;
        end
        th_myfunc_25_9: begin
          th_myfunc_25 <= th_myfunc_25_10;
        end
        th_myfunc_25_10: begin
          $display("Thread %d count = %d", _th_myfunc_25_tid_362, count);
          th_myfunc_25 <= th_myfunc_25_11;
        end
        th_myfunc_25_11: begin
          th_myfunc_25 <= th_myfunc_25_12;
        end
        th_myfunc_25_12: begin
          $display("Thread %d Unlock", _th_myfunc_25_tid_362);
          th_myfunc_25 <= th_myfunc_25_13;
        end
        th_myfunc_25_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 25)) begin
            _th_myfunc_25_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 25)) begin
            th_myfunc_25 <= th_myfunc_25_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_26_1 = 1;
  localparam th_myfunc_26_2 = 2;
  localparam th_myfunc_26_3 = 3;
  localparam th_myfunc_26_4 = 4;
  localparam th_myfunc_26_5 = 5;
  localparam th_myfunc_26_6 = 6;
  localparam th_myfunc_26_7 = 7;
  localparam th_myfunc_26_8 = 8;
  localparam th_myfunc_26_9 = 9;
  localparam th_myfunc_26_10 = 10;
  localparam th_myfunc_26_11 = 11;
  localparam th_myfunc_26_12 = 12;
  localparam th_myfunc_26_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_26 <= th_myfunc_26_init;
      _th_myfunc_26_called <= 0;
      _th_myfunc_26_tid_365 <= 0;
      _th_myfunc_26_tid_366 <= 0;
      _th_myfunc_26_time_367 <= 0;
      _th_myfunc_26_i_368 <= 0;
    end else begin
      case(th_myfunc_26)
        th_myfunc_26_init: begin
          if(_th_myfunc_start[26] && (th_blink == 10)) begin
            _th_myfunc_26_called <= 1;
          end 
          if(_th_myfunc_start[26] && (th_blink == 10)) begin
            _th_myfunc_26_tid_365 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[26]) begin
            th_myfunc_26 <= th_myfunc_26_1;
          end 
        end
        th_myfunc_26_1: begin
          _th_myfunc_26_tid_366 <= _th_myfunc_26_tid_365;
          th_myfunc_26 <= th_myfunc_26_2;
        end
        th_myfunc_26_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 26)) begin
            th_myfunc_26 <= th_myfunc_26_3;
          end 
        end
        th_myfunc_26_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 26))) begin
            th_myfunc_26 <= th_myfunc_26_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 26)) begin
            th_myfunc_26 <= th_myfunc_26_4;
          end 
        end
        th_myfunc_26_4: begin
          $display("Thread %d Lock", _th_myfunc_26_tid_366);
          th_myfunc_26 <= th_myfunc_26_5;
        end
        th_myfunc_26_5: begin
          _th_myfunc_26_time_367 <= sw;
          th_myfunc_26 <= th_myfunc_26_6;
        end
        th_myfunc_26_6: begin
          _th_myfunc_26_i_368 <= 0;
          th_myfunc_26 <= th_myfunc_26_7;
        end
        th_myfunc_26_7: begin
          if(_th_myfunc_26_i_368 < _th_myfunc_26_time_367) begin
            th_myfunc_26 <= th_myfunc_26_8;
          end else begin
            th_myfunc_26 <= th_myfunc_26_9;
          end
        end
        th_myfunc_26_8: begin
          _th_myfunc_26_i_368 <= _th_myfunc_26_i_368 + 1;
          th_myfunc_26 <= th_myfunc_26_7;
        end
        th_myfunc_26_9: begin
          th_myfunc_26 <= th_myfunc_26_10;
        end
        th_myfunc_26_10: begin
          $display("Thread %d count = %d", _th_myfunc_26_tid_366, count);
          th_myfunc_26 <= th_myfunc_26_11;
        end
        th_myfunc_26_11: begin
          th_myfunc_26 <= th_myfunc_26_12;
        end
        th_myfunc_26_12: begin
          $display("Thread %d Unlock", _th_myfunc_26_tid_366);
          th_myfunc_26 <= th_myfunc_26_13;
        end
        th_myfunc_26_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 26)) begin
            _th_myfunc_26_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 26)) begin
            th_myfunc_26 <= th_myfunc_26_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_27_1 = 1;
  localparam th_myfunc_27_2 = 2;
  localparam th_myfunc_27_3 = 3;
  localparam th_myfunc_27_4 = 4;
  localparam th_myfunc_27_5 = 5;
  localparam th_myfunc_27_6 = 6;
  localparam th_myfunc_27_7 = 7;
  localparam th_myfunc_27_8 = 8;
  localparam th_myfunc_27_9 = 9;
  localparam th_myfunc_27_10 = 10;
  localparam th_myfunc_27_11 = 11;
  localparam th_myfunc_27_12 = 12;
  localparam th_myfunc_27_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_27 <= th_myfunc_27_init;
      _th_myfunc_27_called <= 0;
      _th_myfunc_27_tid_369 <= 0;
      _th_myfunc_27_tid_370 <= 0;
      _th_myfunc_27_time_371 <= 0;
      _th_myfunc_27_i_372 <= 0;
    end else begin
      case(th_myfunc_27)
        th_myfunc_27_init: begin
          if(_th_myfunc_start[27] && (th_blink == 10)) begin
            _th_myfunc_27_called <= 1;
          end 
          if(_th_myfunc_start[27] && (th_blink == 10)) begin
            _th_myfunc_27_tid_369 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[27]) begin
            th_myfunc_27 <= th_myfunc_27_1;
          end 
        end
        th_myfunc_27_1: begin
          _th_myfunc_27_tid_370 <= _th_myfunc_27_tid_369;
          th_myfunc_27 <= th_myfunc_27_2;
        end
        th_myfunc_27_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 27)) begin
            th_myfunc_27 <= th_myfunc_27_3;
          end 
        end
        th_myfunc_27_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 27))) begin
            th_myfunc_27 <= th_myfunc_27_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 27)) begin
            th_myfunc_27 <= th_myfunc_27_4;
          end 
        end
        th_myfunc_27_4: begin
          $display("Thread %d Lock", _th_myfunc_27_tid_370);
          th_myfunc_27 <= th_myfunc_27_5;
        end
        th_myfunc_27_5: begin
          _th_myfunc_27_time_371 <= sw;
          th_myfunc_27 <= th_myfunc_27_6;
        end
        th_myfunc_27_6: begin
          _th_myfunc_27_i_372 <= 0;
          th_myfunc_27 <= th_myfunc_27_7;
        end
        th_myfunc_27_7: begin
          if(_th_myfunc_27_i_372 < _th_myfunc_27_time_371) begin
            th_myfunc_27 <= th_myfunc_27_8;
          end else begin
            th_myfunc_27 <= th_myfunc_27_9;
          end
        end
        th_myfunc_27_8: begin
          _th_myfunc_27_i_372 <= _th_myfunc_27_i_372 + 1;
          th_myfunc_27 <= th_myfunc_27_7;
        end
        th_myfunc_27_9: begin
          th_myfunc_27 <= th_myfunc_27_10;
        end
        th_myfunc_27_10: begin
          $display("Thread %d count = %d", _th_myfunc_27_tid_370, count);
          th_myfunc_27 <= th_myfunc_27_11;
        end
        th_myfunc_27_11: begin
          th_myfunc_27 <= th_myfunc_27_12;
        end
        th_myfunc_27_12: begin
          $display("Thread %d Unlock", _th_myfunc_27_tid_370);
          th_myfunc_27 <= th_myfunc_27_13;
        end
        th_myfunc_27_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 27)) begin
            _th_myfunc_27_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 27)) begin
            th_myfunc_27 <= th_myfunc_27_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_28_1 = 1;
  localparam th_myfunc_28_2 = 2;
  localparam th_myfunc_28_3 = 3;
  localparam th_myfunc_28_4 = 4;
  localparam th_myfunc_28_5 = 5;
  localparam th_myfunc_28_6 = 6;
  localparam th_myfunc_28_7 = 7;
  localparam th_myfunc_28_8 = 8;
  localparam th_myfunc_28_9 = 9;
  localparam th_myfunc_28_10 = 10;
  localparam th_myfunc_28_11 = 11;
  localparam th_myfunc_28_12 = 12;
  localparam th_myfunc_28_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_28 <= th_myfunc_28_init;
      _th_myfunc_28_called <= 0;
      _th_myfunc_28_tid_373 <= 0;
      _th_myfunc_28_tid_374 <= 0;
      _th_myfunc_28_time_375 <= 0;
      _th_myfunc_28_i_376 <= 0;
    end else begin
      case(th_myfunc_28)
        th_myfunc_28_init: begin
          if(_th_myfunc_start[28] && (th_blink == 10)) begin
            _th_myfunc_28_called <= 1;
          end 
          if(_th_myfunc_start[28] && (th_blink == 10)) begin
            _th_myfunc_28_tid_373 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[28]) begin
            th_myfunc_28 <= th_myfunc_28_1;
          end 
        end
        th_myfunc_28_1: begin
          _th_myfunc_28_tid_374 <= _th_myfunc_28_tid_373;
          th_myfunc_28 <= th_myfunc_28_2;
        end
        th_myfunc_28_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 28)) begin
            th_myfunc_28 <= th_myfunc_28_3;
          end 
        end
        th_myfunc_28_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 28))) begin
            th_myfunc_28 <= th_myfunc_28_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 28)) begin
            th_myfunc_28 <= th_myfunc_28_4;
          end 
        end
        th_myfunc_28_4: begin
          $display("Thread %d Lock", _th_myfunc_28_tid_374);
          th_myfunc_28 <= th_myfunc_28_5;
        end
        th_myfunc_28_5: begin
          _th_myfunc_28_time_375 <= sw;
          th_myfunc_28 <= th_myfunc_28_6;
        end
        th_myfunc_28_6: begin
          _th_myfunc_28_i_376 <= 0;
          th_myfunc_28 <= th_myfunc_28_7;
        end
        th_myfunc_28_7: begin
          if(_th_myfunc_28_i_376 < _th_myfunc_28_time_375) begin
            th_myfunc_28 <= th_myfunc_28_8;
          end else begin
            th_myfunc_28 <= th_myfunc_28_9;
          end
        end
        th_myfunc_28_8: begin
          _th_myfunc_28_i_376 <= _th_myfunc_28_i_376 + 1;
          th_myfunc_28 <= th_myfunc_28_7;
        end
        th_myfunc_28_9: begin
          th_myfunc_28 <= th_myfunc_28_10;
        end
        th_myfunc_28_10: begin
          $display("Thread %d count = %d", _th_myfunc_28_tid_374, count);
          th_myfunc_28 <= th_myfunc_28_11;
        end
        th_myfunc_28_11: begin
          th_myfunc_28 <= th_myfunc_28_12;
        end
        th_myfunc_28_12: begin
          $display("Thread %d Unlock", _th_myfunc_28_tid_374);
          th_myfunc_28 <= th_myfunc_28_13;
        end
        th_myfunc_28_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 28)) begin
            _th_myfunc_28_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 28)) begin
            th_myfunc_28 <= th_myfunc_28_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_29_1 = 1;
  localparam th_myfunc_29_2 = 2;
  localparam th_myfunc_29_3 = 3;
  localparam th_myfunc_29_4 = 4;
  localparam th_myfunc_29_5 = 5;
  localparam th_myfunc_29_6 = 6;
  localparam th_myfunc_29_7 = 7;
  localparam th_myfunc_29_8 = 8;
  localparam th_myfunc_29_9 = 9;
  localparam th_myfunc_29_10 = 10;
  localparam th_myfunc_29_11 = 11;
  localparam th_myfunc_29_12 = 12;
  localparam th_myfunc_29_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_29 <= th_myfunc_29_init;
      _th_myfunc_29_called <= 0;
      _th_myfunc_29_tid_377 <= 0;
      _th_myfunc_29_tid_378 <= 0;
      _th_myfunc_29_time_379 <= 0;
      _th_myfunc_29_i_380 <= 0;
    end else begin
      case(th_myfunc_29)
        th_myfunc_29_init: begin
          if(_th_myfunc_start[29] && (th_blink == 10)) begin
            _th_myfunc_29_called <= 1;
          end 
          if(_th_myfunc_start[29] && (th_blink == 10)) begin
            _th_myfunc_29_tid_377 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[29]) begin
            th_myfunc_29 <= th_myfunc_29_1;
          end 
        end
        th_myfunc_29_1: begin
          _th_myfunc_29_tid_378 <= _th_myfunc_29_tid_377;
          th_myfunc_29 <= th_myfunc_29_2;
        end
        th_myfunc_29_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 29)) begin
            th_myfunc_29 <= th_myfunc_29_3;
          end 
        end
        th_myfunc_29_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 29))) begin
            th_myfunc_29 <= th_myfunc_29_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 29)) begin
            th_myfunc_29 <= th_myfunc_29_4;
          end 
        end
        th_myfunc_29_4: begin
          $display("Thread %d Lock", _th_myfunc_29_tid_378);
          th_myfunc_29 <= th_myfunc_29_5;
        end
        th_myfunc_29_5: begin
          _th_myfunc_29_time_379 <= sw;
          th_myfunc_29 <= th_myfunc_29_6;
        end
        th_myfunc_29_6: begin
          _th_myfunc_29_i_380 <= 0;
          th_myfunc_29 <= th_myfunc_29_7;
        end
        th_myfunc_29_7: begin
          if(_th_myfunc_29_i_380 < _th_myfunc_29_time_379) begin
            th_myfunc_29 <= th_myfunc_29_8;
          end else begin
            th_myfunc_29 <= th_myfunc_29_9;
          end
        end
        th_myfunc_29_8: begin
          _th_myfunc_29_i_380 <= _th_myfunc_29_i_380 + 1;
          th_myfunc_29 <= th_myfunc_29_7;
        end
        th_myfunc_29_9: begin
          th_myfunc_29 <= th_myfunc_29_10;
        end
        th_myfunc_29_10: begin
          $display("Thread %d count = %d", _th_myfunc_29_tid_378, count);
          th_myfunc_29 <= th_myfunc_29_11;
        end
        th_myfunc_29_11: begin
          th_myfunc_29 <= th_myfunc_29_12;
        end
        th_myfunc_29_12: begin
          $display("Thread %d Unlock", _th_myfunc_29_tid_378);
          th_myfunc_29 <= th_myfunc_29_13;
        end
        th_myfunc_29_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 29)) begin
            _th_myfunc_29_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 29)) begin
            th_myfunc_29 <= th_myfunc_29_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_30_1 = 1;
  localparam th_myfunc_30_2 = 2;
  localparam th_myfunc_30_3 = 3;
  localparam th_myfunc_30_4 = 4;
  localparam th_myfunc_30_5 = 5;
  localparam th_myfunc_30_6 = 6;
  localparam th_myfunc_30_7 = 7;
  localparam th_myfunc_30_8 = 8;
  localparam th_myfunc_30_9 = 9;
  localparam th_myfunc_30_10 = 10;
  localparam th_myfunc_30_11 = 11;
  localparam th_myfunc_30_12 = 12;
  localparam th_myfunc_30_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_30 <= th_myfunc_30_init;
      _th_myfunc_30_called <= 0;
      _th_myfunc_30_tid_381 <= 0;
      _th_myfunc_30_tid_382 <= 0;
      _th_myfunc_30_time_383 <= 0;
      _th_myfunc_30_i_384 <= 0;
    end else begin
      case(th_myfunc_30)
        th_myfunc_30_init: begin
          if(_th_myfunc_start[30] && (th_blink == 10)) begin
            _th_myfunc_30_called <= 1;
          end 
          if(_th_myfunc_start[30] && (th_blink == 10)) begin
            _th_myfunc_30_tid_381 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[30]) begin
            th_myfunc_30 <= th_myfunc_30_1;
          end 
        end
        th_myfunc_30_1: begin
          _th_myfunc_30_tid_382 <= _th_myfunc_30_tid_381;
          th_myfunc_30 <= th_myfunc_30_2;
        end
        th_myfunc_30_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 30)) begin
            th_myfunc_30 <= th_myfunc_30_3;
          end 
        end
        th_myfunc_30_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 30))) begin
            th_myfunc_30 <= th_myfunc_30_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 30)) begin
            th_myfunc_30 <= th_myfunc_30_4;
          end 
        end
        th_myfunc_30_4: begin
          $display("Thread %d Lock", _th_myfunc_30_tid_382);
          th_myfunc_30 <= th_myfunc_30_5;
        end
        th_myfunc_30_5: begin
          _th_myfunc_30_time_383 <= sw;
          th_myfunc_30 <= th_myfunc_30_6;
        end
        th_myfunc_30_6: begin
          _th_myfunc_30_i_384 <= 0;
          th_myfunc_30 <= th_myfunc_30_7;
        end
        th_myfunc_30_7: begin
          if(_th_myfunc_30_i_384 < _th_myfunc_30_time_383) begin
            th_myfunc_30 <= th_myfunc_30_8;
          end else begin
            th_myfunc_30 <= th_myfunc_30_9;
          end
        end
        th_myfunc_30_8: begin
          _th_myfunc_30_i_384 <= _th_myfunc_30_i_384 + 1;
          th_myfunc_30 <= th_myfunc_30_7;
        end
        th_myfunc_30_9: begin
          th_myfunc_30 <= th_myfunc_30_10;
        end
        th_myfunc_30_10: begin
          $display("Thread %d count = %d", _th_myfunc_30_tid_382, count);
          th_myfunc_30 <= th_myfunc_30_11;
        end
        th_myfunc_30_11: begin
          th_myfunc_30 <= th_myfunc_30_12;
        end
        th_myfunc_30_12: begin
          $display("Thread %d Unlock", _th_myfunc_30_tid_382);
          th_myfunc_30 <= th_myfunc_30_13;
        end
        th_myfunc_30_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 30)) begin
            _th_myfunc_30_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 30)) begin
            th_myfunc_30 <= th_myfunc_30_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_31_1 = 1;
  localparam th_myfunc_31_2 = 2;
  localparam th_myfunc_31_3 = 3;
  localparam th_myfunc_31_4 = 4;
  localparam th_myfunc_31_5 = 5;
  localparam th_myfunc_31_6 = 6;
  localparam th_myfunc_31_7 = 7;
  localparam th_myfunc_31_8 = 8;
  localparam th_myfunc_31_9 = 9;
  localparam th_myfunc_31_10 = 10;
  localparam th_myfunc_31_11 = 11;
  localparam th_myfunc_31_12 = 12;
  localparam th_myfunc_31_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_31 <= th_myfunc_31_init;
      _th_myfunc_31_called <= 0;
      _th_myfunc_31_tid_385 <= 0;
      _th_myfunc_31_tid_386 <= 0;
      _th_myfunc_31_time_387 <= 0;
      _th_myfunc_31_i_388 <= 0;
    end else begin
      case(th_myfunc_31)
        th_myfunc_31_init: begin
          if(_th_myfunc_start[31] && (th_blink == 10)) begin
            _th_myfunc_31_called <= 1;
          end 
          if(_th_myfunc_start[31] && (th_blink == 10)) begin
            _th_myfunc_31_tid_385 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[31]) begin
            th_myfunc_31 <= th_myfunc_31_1;
          end 
        end
        th_myfunc_31_1: begin
          _th_myfunc_31_tid_386 <= _th_myfunc_31_tid_385;
          th_myfunc_31 <= th_myfunc_31_2;
        end
        th_myfunc_31_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 31)) begin
            th_myfunc_31 <= th_myfunc_31_3;
          end 
        end
        th_myfunc_31_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 31))) begin
            th_myfunc_31 <= th_myfunc_31_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 31)) begin
            th_myfunc_31 <= th_myfunc_31_4;
          end 
        end
        th_myfunc_31_4: begin
          $display("Thread %d Lock", _th_myfunc_31_tid_386);
          th_myfunc_31 <= th_myfunc_31_5;
        end
        th_myfunc_31_5: begin
          _th_myfunc_31_time_387 <= sw;
          th_myfunc_31 <= th_myfunc_31_6;
        end
        th_myfunc_31_6: begin
          _th_myfunc_31_i_388 <= 0;
          th_myfunc_31 <= th_myfunc_31_7;
        end
        th_myfunc_31_7: begin
          if(_th_myfunc_31_i_388 < _th_myfunc_31_time_387) begin
            th_myfunc_31 <= th_myfunc_31_8;
          end else begin
            th_myfunc_31 <= th_myfunc_31_9;
          end
        end
        th_myfunc_31_8: begin
          _th_myfunc_31_i_388 <= _th_myfunc_31_i_388 + 1;
          th_myfunc_31 <= th_myfunc_31_7;
        end
        th_myfunc_31_9: begin
          th_myfunc_31 <= th_myfunc_31_10;
        end
        th_myfunc_31_10: begin
          $display("Thread %d count = %d", _th_myfunc_31_tid_386, count);
          th_myfunc_31 <= th_myfunc_31_11;
        end
        th_myfunc_31_11: begin
          th_myfunc_31 <= th_myfunc_31_12;
        end
        th_myfunc_31_12: begin
          $display("Thread %d Unlock", _th_myfunc_31_tid_386);
          th_myfunc_31 <= th_myfunc_31_13;
        end
        th_myfunc_31_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 31)) begin
            _th_myfunc_31_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 31)) begin
            th_myfunc_31 <= th_myfunc_31_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_32_1 = 1;
  localparam th_myfunc_32_2 = 2;
  localparam th_myfunc_32_3 = 3;
  localparam th_myfunc_32_4 = 4;
  localparam th_myfunc_32_5 = 5;
  localparam th_myfunc_32_6 = 6;
  localparam th_myfunc_32_7 = 7;
  localparam th_myfunc_32_8 = 8;
  localparam th_myfunc_32_9 = 9;
  localparam th_myfunc_32_10 = 10;
  localparam th_myfunc_32_11 = 11;
  localparam th_myfunc_32_12 = 12;
  localparam th_myfunc_32_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_32 <= th_myfunc_32_init;
      _th_myfunc_32_called <= 0;
      _th_myfunc_32_tid_389 <= 0;
      _th_myfunc_32_tid_390 <= 0;
      _th_myfunc_32_time_391 <= 0;
      _th_myfunc_32_i_392 <= 0;
    end else begin
      case(th_myfunc_32)
        th_myfunc_32_init: begin
          if(_th_myfunc_start[32] && (th_blink == 10)) begin
            _th_myfunc_32_called <= 1;
          end 
          if(_th_myfunc_start[32] && (th_blink == 10)) begin
            _th_myfunc_32_tid_389 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[32]) begin
            th_myfunc_32 <= th_myfunc_32_1;
          end 
        end
        th_myfunc_32_1: begin
          _th_myfunc_32_tid_390 <= _th_myfunc_32_tid_389;
          th_myfunc_32 <= th_myfunc_32_2;
        end
        th_myfunc_32_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 32)) begin
            th_myfunc_32 <= th_myfunc_32_3;
          end 
        end
        th_myfunc_32_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 32))) begin
            th_myfunc_32 <= th_myfunc_32_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 32)) begin
            th_myfunc_32 <= th_myfunc_32_4;
          end 
        end
        th_myfunc_32_4: begin
          $display("Thread %d Lock", _th_myfunc_32_tid_390);
          th_myfunc_32 <= th_myfunc_32_5;
        end
        th_myfunc_32_5: begin
          _th_myfunc_32_time_391 <= sw;
          th_myfunc_32 <= th_myfunc_32_6;
        end
        th_myfunc_32_6: begin
          _th_myfunc_32_i_392 <= 0;
          th_myfunc_32 <= th_myfunc_32_7;
        end
        th_myfunc_32_7: begin
          if(_th_myfunc_32_i_392 < _th_myfunc_32_time_391) begin
            th_myfunc_32 <= th_myfunc_32_8;
          end else begin
            th_myfunc_32 <= th_myfunc_32_9;
          end
        end
        th_myfunc_32_8: begin
          _th_myfunc_32_i_392 <= _th_myfunc_32_i_392 + 1;
          th_myfunc_32 <= th_myfunc_32_7;
        end
        th_myfunc_32_9: begin
          th_myfunc_32 <= th_myfunc_32_10;
        end
        th_myfunc_32_10: begin
          $display("Thread %d count = %d", _th_myfunc_32_tid_390, count);
          th_myfunc_32 <= th_myfunc_32_11;
        end
        th_myfunc_32_11: begin
          th_myfunc_32 <= th_myfunc_32_12;
        end
        th_myfunc_32_12: begin
          $display("Thread %d Unlock", _th_myfunc_32_tid_390);
          th_myfunc_32 <= th_myfunc_32_13;
        end
        th_myfunc_32_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 32)) begin
            _th_myfunc_32_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 32)) begin
            th_myfunc_32 <= th_myfunc_32_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_33_1 = 1;
  localparam th_myfunc_33_2 = 2;
  localparam th_myfunc_33_3 = 3;
  localparam th_myfunc_33_4 = 4;
  localparam th_myfunc_33_5 = 5;
  localparam th_myfunc_33_6 = 6;
  localparam th_myfunc_33_7 = 7;
  localparam th_myfunc_33_8 = 8;
  localparam th_myfunc_33_9 = 9;
  localparam th_myfunc_33_10 = 10;
  localparam th_myfunc_33_11 = 11;
  localparam th_myfunc_33_12 = 12;
  localparam th_myfunc_33_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_33 <= th_myfunc_33_init;
      _th_myfunc_33_called <= 0;
      _th_myfunc_33_tid_393 <= 0;
      _th_myfunc_33_tid_394 <= 0;
      _th_myfunc_33_time_395 <= 0;
      _th_myfunc_33_i_396 <= 0;
    end else begin
      case(th_myfunc_33)
        th_myfunc_33_init: begin
          if(_th_myfunc_start[33] && (th_blink == 10)) begin
            _th_myfunc_33_called <= 1;
          end 
          if(_th_myfunc_start[33] && (th_blink == 10)) begin
            _th_myfunc_33_tid_393 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[33]) begin
            th_myfunc_33 <= th_myfunc_33_1;
          end 
        end
        th_myfunc_33_1: begin
          _th_myfunc_33_tid_394 <= _th_myfunc_33_tid_393;
          th_myfunc_33 <= th_myfunc_33_2;
        end
        th_myfunc_33_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 33)) begin
            th_myfunc_33 <= th_myfunc_33_3;
          end 
        end
        th_myfunc_33_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 33))) begin
            th_myfunc_33 <= th_myfunc_33_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 33)) begin
            th_myfunc_33 <= th_myfunc_33_4;
          end 
        end
        th_myfunc_33_4: begin
          $display("Thread %d Lock", _th_myfunc_33_tid_394);
          th_myfunc_33 <= th_myfunc_33_5;
        end
        th_myfunc_33_5: begin
          _th_myfunc_33_time_395 <= sw;
          th_myfunc_33 <= th_myfunc_33_6;
        end
        th_myfunc_33_6: begin
          _th_myfunc_33_i_396 <= 0;
          th_myfunc_33 <= th_myfunc_33_7;
        end
        th_myfunc_33_7: begin
          if(_th_myfunc_33_i_396 < _th_myfunc_33_time_395) begin
            th_myfunc_33 <= th_myfunc_33_8;
          end else begin
            th_myfunc_33 <= th_myfunc_33_9;
          end
        end
        th_myfunc_33_8: begin
          _th_myfunc_33_i_396 <= _th_myfunc_33_i_396 + 1;
          th_myfunc_33 <= th_myfunc_33_7;
        end
        th_myfunc_33_9: begin
          th_myfunc_33 <= th_myfunc_33_10;
        end
        th_myfunc_33_10: begin
          $display("Thread %d count = %d", _th_myfunc_33_tid_394, count);
          th_myfunc_33 <= th_myfunc_33_11;
        end
        th_myfunc_33_11: begin
          th_myfunc_33 <= th_myfunc_33_12;
        end
        th_myfunc_33_12: begin
          $display("Thread %d Unlock", _th_myfunc_33_tid_394);
          th_myfunc_33 <= th_myfunc_33_13;
        end
        th_myfunc_33_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 33)) begin
            _th_myfunc_33_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 33)) begin
            th_myfunc_33 <= th_myfunc_33_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_34_1 = 1;
  localparam th_myfunc_34_2 = 2;
  localparam th_myfunc_34_3 = 3;
  localparam th_myfunc_34_4 = 4;
  localparam th_myfunc_34_5 = 5;
  localparam th_myfunc_34_6 = 6;
  localparam th_myfunc_34_7 = 7;
  localparam th_myfunc_34_8 = 8;
  localparam th_myfunc_34_9 = 9;
  localparam th_myfunc_34_10 = 10;
  localparam th_myfunc_34_11 = 11;
  localparam th_myfunc_34_12 = 12;
  localparam th_myfunc_34_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_34 <= th_myfunc_34_init;
      _th_myfunc_34_called <= 0;
      _th_myfunc_34_tid_397 <= 0;
      _th_myfunc_34_tid_398 <= 0;
      _th_myfunc_34_time_399 <= 0;
      _th_myfunc_34_i_400 <= 0;
    end else begin
      case(th_myfunc_34)
        th_myfunc_34_init: begin
          if(_th_myfunc_start[34] && (th_blink == 10)) begin
            _th_myfunc_34_called <= 1;
          end 
          if(_th_myfunc_start[34] && (th_blink == 10)) begin
            _th_myfunc_34_tid_397 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[34]) begin
            th_myfunc_34 <= th_myfunc_34_1;
          end 
        end
        th_myfunc_34_1: begin
          _th_myfunc_34_tid_398 <= _th_myfunc_34_tid_397;
          th_myfunc_34 <= th_myfunc_34_2;
        end
        th_myfunc_34_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 34)) begin
            th_myfunc_34 <= th_myfunc_34_3;
          end 
        end
        th_myfunc_34_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 34))) begin
            th_myfunc_34 <= th_myfunc_34_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 34)) begin
            th_myfunc_34 <= th_myfunc_34_4;
          end 
        end
        th_myfunc_34_4: begin
          $display("Thread %d Lock", _th_myfunc_34_tid_398);
          th_myfunc_34 <= th_myfunc_34_5;
        end
        th_myfunc_34_5: begin
          _th_myfunc_34_time_399 <= sw;
          th_myfunc_34 <= th_myfunc_34_6;
        end
        th_myfunc_34_6: begin
          _th_myfunc_34_i_400 <= 0;
          th_myfunc_34 <= th_myfunc_34_7;
        end
        th_myfunc_34_7: begin
          if(_th_myfunc_34_i_400 < _th_myfunc_34_time_399) begin
            th_myfunc_34 <= th_myfunc_34_8;
          end else begin
            th_myfunc_34 <= th_myfunc_34_9;
          end
        end
        th_myfunc_34_8: begin
          _th_myfunc_34_i_400 <= _th_myfunc_34_i_400 + 1;
          th_myfunc_34 <= th_myfunc_34_7;
        end
        th_myfunc_34_9: begin
          th_myfunc_34 <= th_myfunc_34_10;
        end
        th_myfunc_34_10: begin
          $display("Thread %d count = %d", _th_myfunc_34_tid_398, count);
          th_myfunc_34 <= th_myfunc_34_11;
        end
        th_myfunc_34_11: begin
          th_myfunc_34 <= th_myfunc_34_12;
        end
        th_myfunc_34_12: begin
          $display("Thread %d Unlock", _th_myfunc_34_tid_398);
          th_myfunc_34 <= th_myfunc_34_13;
        end
        th_myfunc_34_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 34)) begin
            _th_myfunc_34_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 34)) begin
            th_myfunc_34 <= th_myfunc_34_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_35_1 = 1;
  localparam th_myfunc_35_2 = 2;
  localparam th_myfunc_35_3 = 3;
  localparam th_myfunc_35_4 = 4;
  localparam th_myfunc_35_5 = 5;
  localparam th_myfunc_35_6 = 6;
  localparam th_myfunc_35_7 = 7;
  localparam th_myfunc_35_8 = 8;
  localparam th_myfunc_35_9 = 9;
  localparam th_myfunc_35_10 = 10;
  localparam th_myfunc_35_11 = 11;
  localparam th_myfunc_35_12 = 12;
  localparam th_myfunc_35_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_35 <= th_myfunc_35_init;
      _th_myfunc_35_called <= 0;
      _th_myfunc_35_tid_401 <= 0;
      _th_myfunc_35_tid_402 <= 0;
      _th_myfunc_35_time_403 <= 0;
      _th_myfunc_35_i_404 <= 0;
    end else begin
      case(th_myfunc_35)
        th_myfunc_35_init: begin
          if(_th_myfunc_start[35] && (th_blink == 10)) begin
            _th_myfunc_35_called <= 1;
          end 
          if(_th_myfunc_start[35] && (th_blink == 10)) begin
            _th_myfunc_35_tid_401 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[35]) begin
            th_myfunc_35 <= th_myfunc_35_1;
          end 
        end
        th_myfunc_35_1: begin
          _th_myfunc_35_tid_402 <= _th_myfunc_35_tid_401;
          th_myfunc_35 <= th_myfunc_35_2;
        end
        th_myfunc_35_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 35)) begin
            th_myfunc_35 <= th_myfunc_35_3;
          end 
        end
        th_myfunc_35_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 35))) begin
            th_myfunc_35 <= th_myfunc_35_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 35)) begin
            th_myfunc_35 <= th_myfunc_35_4;
          end 
        end
        th_myfunc_35_4: begin
          $display("Thread %d Lock", _th_myfunc_35_tid_402);
          th_myfunc_35 <= th_myfunc_35_5;
        end
        th_myfunc_35_5: begin
          _th_myfunc_35_time_403 <= sw;
          th_myfunc_35 <= th_myfunc_35_6;
        end
        th_myfunc_35_6: begin
          _th_myfunc_35_i_404 <= 0;
          th_myfunc_35 <= th_myfunc_35_7;
        end
        th_myfunc_35_7: begin
          if(_th_myfunc_35_i_404 < _th_myfunc_35_time_403) begin
            th_myfunc_35 <= th_myfunc_35_8;
          end else begin
            th_myfunc_35 <= th_myfunc_35_9;
          end
        end
        th_myfunc_35_8: begin
          _th_myfunc_35_i_404 <= _th_myfunc_35_i_404 + 1;
          th_myfunc_35 <= th_myfunc_35_7;
        end
        th_myfunc_35_9: begin
          th_myfunc_35 <= th_myfunc_35_10;
        end
        th_myfunc_35_10: begin
          $display("Thread %d count = %d", _th_myfunc_35_tid_402, count);
          th_myfunc_35 <= th_myfunc_35_11;
        end
        th_myfunc_35_11: begin
          th_myfunc_35 <= th_myfunc_35_12;
        end
        th_myfunc_35_12: begin
          $display("Thread %d Unlock", _th_myfunc_35_tid_402);
          th_myfunc_35 <= th_myfunc_35_13;
        end
        th_myfunc_35_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 35)) begin
            _th_myfunc_35_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 35)) begin
            th_myfunc_35 <= th_myfunc_35_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_36_1 = 1;
  localparam th_myfunc_36_2 = 2;
  localparam th_myfunc_36_3 = 3;
  localparam th_myfunc_36_4 = 4;
  localparam th_myfunc_36_5 = 5;
  localparam th_myfunc_36_6 = 6;
  localparam th_myfunc_36_7 = 7;
  localparam th_myfunc_36_8 = 8;
  localparam th_myfunc_36_9 = 9;
  localparam th_myfunc_36_10 = 10;
  localparam th_myfunc_36_11 = 11;
  localparam th_myfunc_36_12 = 12;
  localparam th_myfunc_36_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_36 <= th_myfunc_36_init;
      _th_myfunc_36_called <= 0;
      _th_myfunc_36_tid_405 <= 0;
      _th_myfunc_36_tid_406 <= 0;
      _th_myfunc_36_time_407 <= 0;
      _th_myfunc_36_i_408 <= 0;
    end else begin
      case(th_myfunc_36)
        th_myfunc_36_init: begin
          if(_th_myfunc_start[36] && (th_blink == 10)) begin
            _th_myfunc_36_called <= 1;
          end 
          if(_th_myfunc_start[36] && (th_blink == 10)) begin
            _th_myfunc_36_tid_405 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[36]) begin
            th_myfunc_36 <= th_myfunc_36_1;
          end 
        end
        th_myfunc_36_1: begin
          _th_myfunc_36_tid_406 <= _th_myfunc_36_tid_405;
          th_myfunc_36 <= th_myfunc_36_2;
        end
        th_myfunc_36_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 36)) begin
            th_myfunc_36 <= th_myfunc_36_3;
          end 
        end
        th_myfunc_36_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 36))) begin
            th_myfunc_36 <= th_myfunc_36_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 36)) begin
            th_myfunc_36 <= th_myfunc_36_4;
          end 
        end
        th_myfunc_36_4: begin
          $display("Thread %d Lock", _th_myfunc_36_tid_406);
          th_myfunc_36 <= th_myfunc_36_5;
        end
        th_myfunc_36_5: begin
          _th_myfunc_36_time_407 <= sw;
          th_myfunc_36 <= th_myfunc_36_6;
        end
        th_myfunc_36_6: begin
          _th_myfunc_36_i_408 <= 0;
          th_myfunc_36 <= th_myfunc_36_7;
        end
        th_myfunc_36_7: begin
          if(_th_myfunc_36_i_408 < _th_myfunc_36_time_407) begin
            th_myfunc_36 <= th_myfunc_36_8;
          end else begin
            th_myfunc_36 <= th_myfunc_36_9;
          end
        end
        th_myfunc_36_8: begin
          _th_myfunc_36_i_408 <= _th_myfunc_36_i_408 + 1;
          th_myfunc_36 <= th_myfunc_36_7;
        end
        th_myfunc_36_9: begin
          th_myfunc_36 <= th_myfunc_36_10;
        end
        th_myfunc_36_10: begin
          $display("Thread %d count = %d", _th_myfunc_36_tid_406, count);
          th_myfunc_36 <= th_myfunc_36_11;
        end
        th_myfunc_36_11: begin
          th_myfunc_36 <= th_myfunc_36_12;
        end
        th_myfunc_36_12: begin
          $display("Thread %d Unlock", _th_myfunc_36_tid_406);
          th_myfunc_36 <= th_myfunc_36_13;
        end
        th_myfunc_36_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 36)) begin
            _th_myfunc_36_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 36)) begin
            th_myfunc_36 <= th_myfunc_36_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_37_1 = 1;
  localparam th_myfunc_37_2 = 2;
  localparam th_myfunc_37_3 = 3;
  localparam th_myfunc_37_4 = 4;
  localparam th_myfunc_37_5 = 5;
  localparam th_myfunc_37_6 = 6;
  localparam th_myfunc_37_7 = 7;
  localparam th_myfunc_37_8 = 8;
  localparam th_myfunc_37_9 = 9;
  localparam th_myfunc_37_10 = 10;
  localparam th_myfunc_37_11 = 11;
  localparam th_myfunc_37_12 = 12;
  localparam th_myfunc_37_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_37 <= th_myfunc_37_init;
      _th_myfunc_37_called <= 0;
      _th_myfunc_37_tid_409 <= 0;
      _th_myfunc_37_tid_410 <= 0;
      _th_myfunc_37_time_411 <= 0;
      _th_myfunc_37_i_412 <= 0;
    end else begin
      case(th_myfunc_37)
        th_myfunc_37_init: begin
          if(_th_myfunc_start[37] && (th_blink == 10)) begin
            _th_myfunc_37_called <= 1;
          end 
          if(_th_myfunc_start[37] && (th_blink == 10)) begin
            _th_myfunc_37_tid_409 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[37]) begin
            th_myfunc_37 <= th_myfunc_37_1;
          end 
        end
        th_myfunc_37_1: begin
          _th_myfunc_37_tid_410 <= _th_myfunc_37_tid_409;
          th_myfunc_37 <= th_myfunc_37_2;
        end
        th_myfunc_37_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 37)) begin
            th_myfunc_37 <= th_myfunc_37_3;
          end 
        end
        th_myfunc_37_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 37))) begin
            th_myfunc_37 <= th_myfunc_37_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 37)) begin
            th_myfunc_37 <= th_myfunc_37_4;
          end 
        end
        th_myfunc_37_4: begin
          $display("Thread %d Lock", _th_myfunc_37_tid_410);
          th_myfunc_37 <= th_myfunc_37_5;
        end
        th_myfunc_37_5: begin
          _th_myfunc_37_time_411 <= sw;
          th_myfunc_37 <= th_myfunc_37_6;
        end
        th_myfunc_37_6: begin
          _th_myfunc_37_i_412 <= 0;
          th_myfunc_37 <= th_myfunc_37_7;
        end
        th_myfunc_37_7: begin
          if(_th_myfunc_37_i_412 < _th_myfunc_37_time_411) begin
            th_myfunc_37 <= th_myfunc_37_8;
          end else begin
            th_myfunc_37 <= th_myfunc_37_9;
          end
        end
        th_myfunc_37_8: begin
          _th_myfunc_37_i_412 <= _th_myfunc_37_i_412 + 1;
          th_myfunc_37 <= th_myfunc_37_7;
        end
        th_myfunc_37_9: begin
          th_myfunc_37 <= th_myfunc_37_10;
        end
        th_myfunc_37_10: begin
          $display("Thread %d count = %d", _th_myfunc_37_tid_410, count);
          th_myfunc_37 <= th_myfunc_37_11;
        end
        th_myfunc_37_11: begin
          th_myfunc_37 <= th_myfunc_37_12;
        end
        th_myfunc_37_12: begin
          $display("Thread %d Unlock", _th_myfunc_37_tid_410);
          th_myfunc_37 <= th_myfunc_37_13;
        end
        th_myfunc_37_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 37)) begin
            _th_myfunc_37_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 37)) begin
            th_myfunc_37 <= th_myfunc_37_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_38_1 = 1;
  localparam th_myfunc_38_2 = 2;
  localparam th_myfunc_38_3 = 3;
  localparam th_myfunc_38_4 = 4;
  localparam th_myfunc_38_5 = 5;
  localparam th_myfunc_38_6 = 6;
  localparam th_myfunc_38_7 = 7;
  localparam th_myfunc_38_8 = 8;
  localparam th_myfunc_38_9 = 9;
  localparam th_myfunc_38_10 = 10;
  localparam th_myfunc_38_11 = 11;
  localparam th_myfunc_38_12 = 12;
  localparam th_myfunc_38_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_38 <= th_myfunc_38_init;
      _th_myfunc_38_called <= 0;
      _th_myfunc_38_tid_413 <= 0;
      _th_myfunc_38_tid_414 <= 0;
      _th_myfunc_38_time_415 <= 0;
      _th_myfunc_38_i_416 <= 0;
    end else begin
      case(th_myfunc_38)
        th_myfunc_38_init: begin
          if(_th_myfunc_start[38] && (th_blink == 10)) begin
            _th_myfunc_38_called <= 1;
          end 
          if(_th_myfunc_start[38] && (th_blink == 10)) begin
            _th_myfunc_38_tid_413 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[38]) begin
            th_myfunc_38 <= th_myfunc_38_1;
          end 
        end
        th_myfunc_38_1: begin
          _th_myfunc_38_tid_414 <= _th_myfunc_38_tid_413;
          th_myfunc_38 <= th_myfunc_38_2;
        end
        th_myfunc_38_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 38)) begin
            th_myfunc_38 <= th_myfunc_38_3;
          end 
        end
        th_myfunc_38_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 38))) begin
            th_myfunc_38 <= th_myfunc_38_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 38)) begin
            th_myfunc_38 <= th_myfunc_38_4;
          end 
        end
        th_myfunc_38_4: begin
          $display("Thread %d Lock", _th_myfunc_38_tid_414);
          th_myfunc_38 <= th_myfunc_38_5;
        end
        th_myfunc_38_5: begin
          _th_myfunc_38_time_415 <= sw;
          th_myfunc_38 <= th_myfunc_38_6;
        end
        th_myfunc_38_6: begin
          _th_myfunc_38_i_416 <= 0;
          th_myfunc_38 <= th_myfunc_38_7;
        end
        th_myfunc_38_7: begin
          if(_th_myfunc_38_i_416 < _th_myfunc_38_time_415) begin
            th_myfunc_38 <= th_myfunc_38_8;
          end else begin
            th_myfunc_38 <= th_myfunc_38_9;
          end
        end
        th_myfunc_38_8: begin
          _th_myfunc_38_i_416 <= _th_myfunc_38_i_416 + 1;
          th_myfunc_38 <= th_myfunc_38_7;
        end
        th_myfunc_38_9: begin
          th_myfunc_38 <= th_myfunc_38_10;
        end
        th_myfunc_38_10: begin
          $display("Thread %d count = %d", _th_myfunc_38_tid_414, count);
          th_myfunc_38 <= th_myfunc_38_11;
        end
        th_myfunc_38_11: begin
          th_myfunc_38 <= th_myfunc_38_12;
        end
        th_myfunc_38_12: begin
          $display("Thread %d Unlock", _th_myfunc_38_tid_414);
          th_myfunc_38 <= th_myfunc_38_13;
        end
        th_myfunc_38_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 38)) begin
            _th_myfunc_38_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 38)) begin
            th_myfunc_38 <= th_myfunc_38_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_39_1 = 1;
  localparam th_myfunc_39_2 = 2;
  localparam th_myfunc_39_3 = 3;
  localparam th_myfunc_39_4 = 4;
  localparam th_myfunc_39_5 = 5;
  localparam th_myfunc_39_6 = 6;
  localparam th_myfunc_39_7 = 7;
  localparam th_myfunc_39_8 = 8;
  localparam th_myfunc_39_9 = 9;
  localparam th_myfunc_39_10 = 10;
  localparam th_myfunc_39_11 = 11;
  localparam th_myfunc_39_12 = 12;
  localparam th_myfunc_39_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_39 <= th_myfunc_39_init;
      _th_myfunc_39_called <= 0;
      _th_myfunc_39_tid_417 <= 0;
      _th_myfunc_39_tid_418 <= 0;
      _th_myfunc_39_time_419 <= 0;
      _th_myfunc_39_i_420 <= 0;
    end else begin
      case(th_myfunc_39)
        th_myfunc_39_init: begin
          if(_th_myfunc_start[39] && (th_blink == 10)) begin
            _th_myfunc_39_called <= 1;
          end 
          if(_th_myfunc_start[39] && (th_blink == 10)) begin
            _th_myfunc_39_tid_417 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[39]) begin
            th_myfunc_39 <= th_myfunc_39_1;
          end 
        end
        th_myfunc_39_1: begin
          _th_myfunc_39_tid_418 <= _th_myfunc_39_tid_417;
          th_myfunc_39 <= th_myfunc_39_2;
        end
        th_myfunc_39_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 39)) begin
            th_myfunc_39 <= th_myfunc_39_3;
          end 
        end
        th_myfunc_39_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 39))) begin
            th_myfunc_39 <= th_myfunc_39_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 39)) begin
            th_myfunc_39 <= th_myfunc_39_4;
          end 
        end
        th_myfunc_39_4: begin
          $display("Thread %d Lock", _th_myfunc_39_tid_418);
          th_myfunc_39 <= th_myfunc_39_5;
        end
        th_myfunc_39_5: begin
          _th_myfunc_39_time_419 <= sw;
          th_myfunc_39 <= th_myfunc_39_6;
        end
        th_myfunc_39_6: begin
          _th_myfunc_39_i_420 <= 0;
          th_myfunc_39 <= th_myfunc_39_7;
        end
        th_myfunc_39_7: begin
          if(_th_myfunc_39_i_420 < _th_myfunc_39_time_419) begin
            th_myfunc_39 <= th_myfunc_39_8;
          end else begin
            th_myfunc_39 <= th_myfunc_39_9;
          end
        end
        th_myfunc_39_8: begin
          _th_myfunc_39_i_420 <= _th_myfunc_39_i_420 + 1;
          th_myfunc_39 <= th_myfunc_39_7;
        end
        th_myfunc_39_9: begin
          th_myfunc_39 <= th_myfunc_39_10;
        end
        th_myfunc_39_10: begin
          $display("Thread %d count = %d", _th_myfunc_39_tid_418, count);
          th_myfunc_39 <= th_myfunc_39_11;
        end
        th_myfunc_39_11: begin
          th_myfunc_39 <= th_myfunc_39_12;
        end
        th_myfunc_39_12: begin
          $display("Thread %d Unlock", _th_myfunc_39_tid_418);
          th_myfunc_39 <= th_myfunc_39_13;
        end
        th_myfunc_39_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 39)) begin
            _th_myfunc_39_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 39)) begin
            th_myfunc_39 <= th_myfunc_39_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_40_1 = 1;
  localparam th_myfunc_40_2 = 2;
  localparam th_myfunc_40_3 = 3;
  localparam th_myfunc_40_4 = 4;
  localparam th_myfunc_40_5 = 5;
  localparam th_myfunc_40_6 = 6;
  localparam th_myfunc_40_7 = 7;
  localparam th_myfunc_40_8 = 8;
  localparam th_myfunc_40_9 = 9;
  localparam th_myfunc_40_10 = 10;
  localparam th_myfunc_40_11 = 11;
  localparam th_myfunc_40_12 = 12;
  localparam th_myfunc_40_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_40 <= th_myfunc_40_init;
      _th_myfunc_40_called <= 0;
      _th_myfunc_40_tid_421 <= 0;
      _th_myfunc_40_tid_422 <= 0;
      _th_myfunc_40_time_423 <= 0;
      _th_myfunc_40_i_424 <= 0;
    end else begin
      case(th_myfunc_40)
        th_myfunc_40_init: begin
          if(_th_myfunc_start[40] && (th_blink == 10)) begin
            _th_myfunc_40_called <= 1;
          end 
          if(_th_myfunc_start[40] && (th_blink == 10)) begin
            _th_myfunc_40_tid_421 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[40]) begin
            th_myfunc_40 <= th_myfunc_40_1;
          end 
        end
        th_myfunc_40_1: begin
          _th_myfunc_40_tid_422 <= _th_myfunc_40_tid_421;
          th_myfunc_40 <= th_myfunc_40_2;
        end
        th_myfunc_40_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 40)) begin
            th_myfunc_40 <= th_myfunc_40_3;
          end 
        end
        th_myfunc_40_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 40))) begin
            th_myfunc_40 <= th_myfunc_40_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 40)) begin
            th_myfunc_40 <= th_myfunc_40_4;
          end 
        end
        th_myfunc_40_4: begin
          $display("Thread %d Lock", _th_myfunc_40_tid_422);
          th_myfunc_40 <= th_myfunc_40_5;
        end
        th_myfunc_40_5: begin
          _th_myfunc_40_time_423 <= sw;
          th_myfunc_40 <= th_myfunc_40_6;
        end
        th_myfunc_40_6: begin
          _th_myfunc_40_i_424 <= 0;
          th_myfunc_40 <= th_myfunc_40_7;
        end
        th_myfunc_40_7: begin
          if(_th_myfunc_40_i_424 < _th_myfunc_40_time_423) begin
            th_myfunc_40 <= th_myfunc_40_8;
          end else begin
            th_myfunc_40 <= th_myfunc_40_9;
          end
        end
        th_myfunc_40_8: begin
          _th_myfunc_40_i_424 <= _th_myfunc_40_i_424 + 1;
          th_myfunc_40 <= th_myfunc_40_7;
        end
        th_myfunc_40_9: begin
          th_myfunc_40 <= th_myfunc_40_10;
        end
        th_myfunc_40_10: begin
          $display("Thread %d count = %d", _th_myfunc_40_tid_422, count);
          th_myfunc_40 <= th_myfunc_40_11;
        end
        th_myfunc_40_11: begin
          th_myfunc_40 <= th_myfunc_40_12;
        end
        th_myfunc_40_12: begin
          $display("Thread %d Unlock", _th_myfunc_40_tid_422);
          th_myfunc_40 <= th_myfunc_40_13;
        end
        th_myfunc_40_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 40)) begin
            _th_myfunc_40_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 40)) begin
            th_myfunc_40 <= th_myfunc_40_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_41_1 = 1;
  localparam th_myfunc_41_2 = 2;
  localparam th_myfunc_41_3 = 3;
  localparam th_myfunc_41_4 = 4;
  localparam th_myfunc_41_5 = 5;
  localparam th_myfunc_41_6 = 6;
  localparam th_myfunc_41_7 = 7;
  localparam th_myfunc_41_8 = 8;
  localparam th_myfunc_41_9 = 9;
  localparam th_myfunc_41_10 = 10;
  localparam th_myfunc_41_11 = 11;
  localparam th_myfunc_41_12 = 12;
  localparam th_myfunc_41_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_41 <= th_myfunc_41_init;
      _th_myfunc_41_called <= 0;
      _th_myfunc_41_tid_425 <= 0;
      _th_myfunc_41_tid_426 <= 0;
      _th_myfunc_41_time_427 <= 0;
      _th_myfunc_41_i_428 <= 0;
    end else begin
      case(th_myfunc_41)
        th_myfunc_41_init: begin
          if(_th_myfunc_start[41] && (th_blink == 10)) begin
            _th_myfunc_41_called <= 1;
          end 
          if(_th_myfunc_start[41] && (th_blink == 10)) begin
            _th_myfunc_41_tid_425 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[41]) begin
            th_myfunc_41 <= th_myfunc_41_1;
          end 
        end
        th_myfunc_41_1: begin
          _th_myfunc_41_tid_426 <= _th_myfunc_41_tid_425;
          th_myfunc_41 <= th_myfunc_41_2;
        end
        th_myfunc_41_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 41)) begin
            th_myfunc_41 <= th_myfunc_41_3;
          end 
        end
        th_myfunc_41_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 41))) begin
            th_myfunc_41 <= th_myfunc_41_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 41)) begin
            th_myfunc_41 <= th_myfunc_41_4;
          end 
        end
        th_myfunc_41_4: begin
          $display("Thread %d Lock", _th_myfunc_41_tid_426);
          th_myfunc_41 <= th_myfunc_41_5;
        end
        th_myfunc_41_5: begin
          _th_myfunc_41_time_427 <= sw;
          th_myfunc_41 <= th_myfunc_41_6;
        end
        th_myfunc_41_6: begin
          _th_myfunc_41_i_428 <= 0;
          th_myfunc_41 <= th_myfunc_41_7;
        end
        th_myfunc_41_7: begin
          if(_th_myfunc_41_i_428 < _th_myfunc_41_time_427) begin
            th_myfunc_41 <= th_myfunc_41_8;
          end else begin
            th_myfunc_41 <= th_myfunc_41_9;
          end
        end
        th_myfunc_41_8: begin
          _th_myfunc_41_i_428 <= _th_myfunc_41_i_428 + 1;
          th_myfunc_41 <= th_myfunc_41_7;
        end
        th_myfunc_41_9: begin
          th_myfunc_41 <= th_myfunc_41_10;
        end
        th_myfunc_41_10: begin
          $display("Thread %d count = %d", _th_myfunc_41_tid_426, count);
          th_myfunc_41 <= th_myfunc_41_11;
        end
        th_myfunc_41_11: begin
          th_myfunc_41 <= th_myfunc_41_12;
        end
        th_myfunc_41_12: begin
          $display("Thread %d Unlock", _th_myfunc_41_tid_426);
          th_myfunc_41 <= th_myfunc_41_13;
        end
        th_myfunc_41_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 41)) begin
            _th_myfunc_41_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 41)) begin
            th_myfunc_41 <= th_myfunc_41_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_42_1 = 1;
  localparam th_myfunc_42_2 = 2;
  localparam th_myfunc_42_3 = 3;
  localparam th_myfunc_42_4 = 4;
  localparam th_myfunc_42_5 = 5;
  localparam th_myfunc_42_6 = 6;
  localparam th_myfunc_42_7 = 7;
  localparam th_myfunc_42_8 = 8;
  localparam th_myfunc_42_9 = 9;
  localparam th_myfunc_42_10 = 10;
  localparam th_myfunc_42_11 = 11;
  localparam th_myfunc_42_12 = 12;
  localparam th_myfunc_42_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_42 <= th_myfunc_42_init;
      _th_myfunc_42_called <= 0;
      _th_myfunc_42_tid_429 <= 0;
      _th_myfunc_42_tid_430 <= 0;
      _th_myfunc_42_time_431 <= 0;
      _th_myfunc_42_i_432 <= 0;
    end else begin
      case(th_myfunc_42)
        th_myfunc_42_init: begin
          if(_th_myfunc_start[42] && (th_blink == 10)) begin
            _th_myfunc_42_called <= 1;
          end 
          if(_th_myfunc_start[42] && (th_blink == 10)) begin
            _th_myfunc_42_tid_429 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[42]) begin
            th_myfunc_42 <= th_myfunc_42_1;
          end 
        end
        th_myfunc_42_1: begin
          _th_myfunc_42_tid_430 <= _th_myfunc_42_tid_429;
          th_myfunc_42 <= th_myfunc_42_2;
        end
        th_myfunc_42_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 42)) begin
            th_myfunc_42 <= th_myfunc_42_3;
          end 
        end
        th_myfunc_42_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 42))) begin
            th_myfunc_42 <= th_myfunc_42_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 42)) begin
            th_myfunc_42 <= th_myfunc_42_4;
          end 
        end
        th_myfunc_42_4: begin
          $display("Thread %d Lock", _th_myfunc_42_tid_430);
          th_myfunc_42 <= th_myfunc_42_5;
        end
        th_myfunc_42_5: begin
          _th_myfunc_42_time_431 <= sw;
          th_myfunc_42 <= th_myfunc_42_6;
        end
        th_myfunc_42_6: begin
          _th_myfunc_42_i_432 <= 0;
          th_myfunc_42 <= th_myfunc_42_7;
        end
        th_myfunc_42_7: begin
          if(_th_myfunc_42_i_432 < _th_myfunc_42_time_431) begin
            th_myfunc_42 <= th_myfunc_42_8;
          end else begin
            th_myfunc_42 <= th_myfunc_42_9;
          end
        end
        th_myfunc_42_8: begin
          _th_myfunc_42_i_432 <= _th_myfunc_42_i_432 + 1;
          th_myfunc_42 <= th_myfunc_42_7;
        end
        th_myfunc_42_9: begin
          th_myfunc_42 <= th_myfunc_42_10;
        end
        th_myfunc_42_10: begin
          $display("Thread %d count = %d", _th_myfunc_42_tid_430, count);
          th_myfunc_42 <= th_myfunc_42_11;
        end
        th_myfunc_42_11: begin
          th_myfunc_42 <= th_myfunc_42_12;
        end
        th_myfunc_42_12: begin
          $display("Thread %d Unlock", _th_myfunc_42_tid_430);
          th_myfunc_42 <= th_myfunc_42_13;
        end
        th_myfunc_42_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 42)) begin
            _th_myfunc_42_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 42)) begin
            th_myfunc_42 <= th_myfunc_42_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_43_1 = 1;
  localparam th_myfunc_43_2 = 2;
  localparam th_myfunc_43_3 = 3;
  localparam th_myfunc_43_4 = 4;
  localparam th_myfunc_43_5 = 5;
  localparam th_myfunc_43_6 = 6;
  localparam th_myfunc_43_7 = 7;
  localparam th_myfunc_43_8 = 8;
  localparam th_myfunc_43_9 = 9;
  localparam th_myfunc_43_10 = 10;
  localparam th_myfunc_43_11 = 11;
  localparam th_myfunc_43_12 = 12;
  localparam th_myfunc_43_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_43 <= th_myfunc_43_init;
      _th_myfunc_43_called <= 0;
      _th_myfunc_43_tid_433 <= 0;
      _th_myfunc_43_tid_434 <= 0;
      _th_myfunc_43_time_435 <= 0;
      _th_myfunc_43_i_436 <= 0;
    end else begin
      case(th_myfunc_43)
        th_myfunc_43_init: begin
          if(_th_myfunc_start[43] && (th_blink == 10)) begin
            _th_myfunc_43_called <= 1;
          end 
          if(_th_myfunc_start[43] && (th_blink == 10)) begin
            _th_myfunc_43_tid_433 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[43]) begin
            th_myfunc_43 <= th_myfunc_43_1;
          end 
        end
        th_myfunc_43_1: begin
          _th_myfunc_43_tid_434 <= _th_myfunc_43_tid_433;
          th_myfunc_43 <= th_myfunc_43_2;
        end
        th_myfunc_43_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 43)) begin
            th_myfunc_43 <= th_myfunc_43_3;
          end 
        end
        th_myfunc_43_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 43))) begin
            th_myfunc_43 <= th_myfunc_43_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 43)) begin
            th_myfunc_43 <= th_myfunc_43_4;
          end 
        end
        th_myfunc_43_4: begin
          $display("Thread %d Lock", _th_myfunc_43_tid_434);
          th_myfunc_43 <= th_myfunc_43_5;
        end
        th_myfunc_43_5: begin
          _th_myfunc_43_time_435 <= sw;
          th_myfunc_43 <= th_myfunc_43_6;
        end
        th_myfunc_43_6: begin
          _th_myfunc_43_i_436 <= 0;
          th_myfunc_43 <= th_myfunc_43_7;
        end
        th_myfunc_43_7: begin
          if(_th_myfunc_43_i_436 < _th_myfunc_43_time_435) begin
            th_myfunc_43 <= th_myfunc_43_8;
          end else begin
            th_myfunc_43 <= th_myfunc_43_9;
          end
        end
        th_myfunc_43_8: begin
          _th_myfunc_43_i_436 <= _th_myfunc_43_i_436 + 1;
          th_myfunc_43 <= th_myfunc_43_7;
        end
        th_myfunc_43_9: begin
          th_myfunc_43 <= th_myfunc_43_10;
        end
        th_myfunc_43_10: begin
          $display("Thread %d count = %d", _th_myfunc_43_tid_434, count);
          th_myfunc_43 <= th_myfunc_43_11;
        end
        th_myfunc_43_11: begin
          th_myfunc_43 <= th_myfunc_43_12;
        end
        th_myfunc_43_12: begin
          $display("Thread %d Unlock", _th_myfunc_43_tid_434);
          th_myfunc_43 <= th_myfunc_43_13;
        end
        th_myfunc_43_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 43)) begin
            _th_myfunc_43_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 43)) begin
            th_myfunc_43 <= th_myfunc_43_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_44_1 = 1;
  localparam th_myfunc_44_2 = 2;
  localparam th_myfunc_44_3 = 3;
  localparam th_myfunc_44_4 = 4;
  localparam th_myfunc_44_5 = 5;
  localparam th_myfunc_44_6 = 6;
  localparam th_myfunc_44_7 = 7;
  localparam th_myfunc_44_8 = 8;
  localparam th_myfunc_44_9 = 9;
  localparam th_myfunc_44_10 = 10;
  localparam th_myfunc_44_11 = 11;
  localparam th_myfunc_44_12 = 12;
  localparam th_myfunc_44_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_44 <= th_myfunc_44_init;
      _th_myfunc_44_called <= 0;
      _th_myfunc_44_tid_437 <= 0;
      _th_myfunc_44_tid_438 <= 0;
      _th_myfunc_44_time_439 <= 0;
      _th_myfunc_44_i_440 <= 0;
    end else begin
      case(th_myfunc_44)
        th_myfunc_44_init: begin
          if(_th_myfunc_start[44] && (th_blink == 10)) begin
            _th_myfunc_44_called <= 1;
          end 
          if(_th_myfunc_start[44] && (th_blink == 10)) begin
            _th_myfunc_44_tid_437 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[44]) begin
            th_myfunc_44 <= th_myfunc_44_1;
          end 
        end
        th_myfunc_44_1: begin
          _th_myfunc_44_tid_438 <= _th_myfunc_44_tid_437;
          th_myfunc_44 <= th_myfunc_44_2;
        end
        th_myfunc_44_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 44)) begin
            th_myfunc_44 <= th_myfunc_44_3;
          end 
        end
        th_myfunc_44_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 44))) begin
            th_myfunc_44 <= th_myfunc_44_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 44)) begin
            th_myfunc_44 <= th_myfunc_44_4;
          end 
        end
        th_myfunc_44_4: begin
          $display("Thread %d Lock", _th_myfunc_44_tid_438);
          th_myfunc_44 <= th_myfunc_44_5;
        end
        th_myfunc_44_5: begin
          _th_myfunc_44_time_439 <= sw;
          th_myfunc_44 <= th_myfunc_44_6;
        end
        th_myfunc_44_6: begin
          _th_myfunc_44_i_440 <= 0;
          th_myfunc_44 <= th_myfunc_44_7;
        end
        th_myfunc_44_7: begin
          if(_th_myfunc_44_i_440 < _th_myfunc_44_time_439) begin
            th_myfunc_44 <= th_myfunc_44_8;
          end else begin
            th_myfunc_44 <= th_myfunc_44_9;
          end
        end
        th_myfunc_44_8: begin
          _th_myfunc_44_i_440 <= _th_myfunc_44_i_440 + 1;
          th_myfunc_44 <= th_myfunc_44_7;
        end
        th_myfunc_44_9: begin
          th_myfunc_44 <= th_myfunc_44_10;
        end
        th_myfunc_44_10: begin
          $display("Thread %d count = %d", _th_myfunc_44_tid_438, count);
          th_myfunc_44 <= th_myfunc_44_11;
        end
        th_myfunc_44_11: begin
          th_myfunc_44 <= th_myfunc_44_12;
        end
        th_myfunc_44_12: begin
          $display("Thread %d Unlock", _th_myfunc_44_tid_438);
          th_myfunc_44 <= th_myfunc_44_13;
        end
        th_myfunc_44_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 44)) begin
            _th_myfunc_44_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 44)) begin
            th_myfunc_44 <= th_myfunc_44_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_45_1 = 1;
  localparam th_myfunc_45_2 = 2;
  localparam th_myfunc_45_3 = 3;
  localparam th_myfunc_45_4 = 4;
  localparam th_myfunc_45_5 = 5;
  localparam th_myfunc_45_6 = 6;
  localparam th_myfunc_45_7 = 7;
  localparam th_myfunc_45_8 = 8;
  localparam th_myfunc_45_9 = 9;
  localparam th_myfunc_45_10 = 10;
  localparam th_myfunc_45_11 = 11;
  localparam th_myfunc_45_12 = 12;
  localparam th_myfunc_45_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_45 <= th_myfunc_45_init;
      _th_myfunc_45_called <= 0;
      _th_myfunc_45_tid_441 <= 0;
      _th_myfunc_45_tid_442 <= 0;
      _th_myfunc_45_time_443 <= 0;
      _th_myfunc_45_i_444 <= 0;
    end else begin
      case(th_myfunc_45)
        th_myfunc_45_init: begin
          if(_th_myfunc_start[45] && (th_blink == 10)) begin
            _th_myfunc_45_called <= 1;
          end 
          if(_th_myfunc_start[45] && (th_blink == 10)) begin
            _th_myfunc_45_tid_441 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[45]) begin
            th_myfunc_45 <= th_myfunc_45_1;
          end 
        end
        th_myfunc_45_1: begin
          _th_myfunc_45_tid_442 <= _th_myfunc_45_tid_441;
          th_myfunc_45 <= th_myfunc_45_2;
        end
        th_myfunc_45_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 45)) begin
            th_myfunc_45 <= th_myfunc_45_3;
          end 
        end
        th_myfunc_45_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 45))) begin
            th_myfunc_45 <= th_myfunc_45_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 45)) begin
            th_myfunc_45 <= th_myfunc_45_4;
          end 
        end
        th_myfunc_45_4: begin
          $display("Thread %d Lock", _th_myfunc_45_tid_442);
          th_myfunc_45 <= th_myfunc_45_5;
        end
        th_myfunc_45_5: begin
          _th_myfunc_45_time_443 <= sw;
          th_myfunc_45 <= th_myfunc_45_6;
        end
        th_myfunc_45_6: begin
          _th_myfunc_45_i_444 <= 0;
          th_myfunc_45 <= th_myfunc_45_7;
        end
        th_myfunc_45_7: begin
          if(_th_myfunc_45_i_444 < _th_myfunc_45_time_443) begin
            th_myfunc_45 <= th_myfunc_45_8;
          end else begin
            th_myfunc_45 <= th_myfunc_45_9;
          end
        end
        th_myfunc_45_8: begin
          _th_myfunc_45_i_444 <= _th_myfunc_45_i_444 + 1;
          th_myfunc_45 <= th_myfunc_45_7;
        end
        th_myfunc_45_9: begin
          th_myfunc_45 <= th_myfunc_45_10;
        end
        th_myfunc_45_10: begin
          $display("Thread %d count = %d", _th_myfunc_45_tid_442, count);
          th_myfunc_45 <= th_myfunc_45_11;
        end
        th_myfunc_45_11: begin
          th_myfunc_45 <= th_myfunc_45_12;
        end
        th_myfunc_45_12: begin
          $display("Thread %d Unlock", _th_myfunc_45_tid_442);
          th_myfunc_45 <= th_myfunc_45_13;
        end
        th_myfunc_45_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 45)) begin
            _th_myfunc_45_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 45)) begin
            th_myfunc_45 <= th_myfunc_45_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_46_1 = 1;
  localparam th_myfunc_46_2 = 2;
  localparam th_myfunc_46_3 = 3;
  localparam th_myfunc_46_4 = 4;
  localparam th_myfunc_46_5 = 5;
  localparam th_myfunc_46_6 = 6;
  localparam th_myfunc_46_7 = 7;
  localparam th_myfunc_46_8 = 8;
  localparam th_myfunc_46_9 = 9;
  localparam th_myfunc_46_10 = 10;
  localparam th_myfunc_46_11 = 11;
  localparam th_myfunc_46_12 = 12;
  localparam th_myfunc_46_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_46 <= th_myfunc_46_init;
      _th_myfunc_46_called <= 0;
      _th_myfunc_46_tid_445 <= 0;
      _th_myfunc_46_tid_446 <= 0;
      _th_myfunc_46_time_447 <= 0;
      _th_myfunc_46_i_448 <= 0;
    end else begin
      case(th_myfunc_46)
        th_myfunc_46_init: begin
          if(_th_myfunc_start[46] && (th_blink == 10)) begin
            _th_myfunc_46_called <= 1;
          end 
          if(_th_myfunc_start[46] && (th_blink == 10)) begin
            _th_myfunc_46_tid_445 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[46]) begin
            th_myfunc_46 <= th_myfunc_46_1;
          end 
        end
        th_myfunc_46_1: begin
          _th_myfunc_46_tid_446 <= _th_myfunc_46_tid_445;
          th_myfunc_46 <= th_myfunc_46_2;
        end
        th_myfunc_46_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 46)) begin
            th_myfunc_46 <= th_myfunc_46_3;
          end 
        end
        th_myfunc_46_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 46))) begin
            th_myfunc_46 <= th_myfunc_46_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 46)) begin
            th_myfunc_46 <= th_myfunc_46_4;
          end 
        end
        th_myfunc_46_4: begin
          $display("Thread %d Lock", _th_myfunc_46_tid_446);
          th_myfunc_46 <= th_myfunc_46_5;
        end
        th_myfunc_46_5: begin
          _th_myfunc_46_time_447 <= sw;
          th_myfunc_46 <= th_myfunc_46_6;
        end
        th_myfunc_46_6: begin
          _th_myfunc_46_i_448 <= 0;
          th_myfunc_46 <= th_myfunc_46_7;
        end
        th_myfunc_46_7: begin
          if(_th_myfunc_46_i_448 < _th_myfunc_46_time_447) begin
            th_myfunc_46 <= th_myfunc_46_8;
          end else begin
            th_myfunc_46 <= th_myfunc_46_9;
          end
        end
        th_myfunc_46_8: begin
          _th_myfunc_46_i_448 <= _th_myfunc_46_i_448 + 1;
          th_myfunc_46 <= th_myfunc_46_7;
        end
        th_myfunc_46_9: begin
          th_myfunc_46 <= th_myfunc_46_10;
        end
        th_myfunc_46_10: begin
          $display("Thread %d count = %d", _th_myfunc_46_tid_446, count);
          th_myfunc_46 <= th_myfunc_46_11;
        end
        th_myfunc_46_11: begin
          th_myfunc_46 <= th_myfunc_46_12;
        end
        th_myfunc_46_12: begin
          $display("Thread %d Unlock", _th_myfunc_46_tid_446);
          th_myfunc_46 <= th_myfunc_46_13;
        end
        th_myfunc_46_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 46)) begin
            _th_myfunc_46_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 46)) begin
            th_myfunc_46 <= th_myfunc_46_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_47_1 = 1;
  localparam th_myfunc_47_2 = 2;
  localparam th_myfunc_47_3 = 3;
  localparam th_myfunc_47_4 = 4;
  localparam th_myfunc_47_5 = 5;
  localparam th_myfunc_47_6 = 6;
  localparam th_myfunc_47_7 = 7;
  localparam th_myfunc_47_8 = 8;
  localparam th_myfunc_47_9 = 9;
  localparam th_myfunc_47_10 = 10;
  localparam th_myfunc_47_11 = 11;
  localparam th_myfunc_47_12 = 12;
  localparam th_myfunc_47_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_47 <= th_myfunc_47_init;
      _th_myfunc_47_called <= 0;
      _th_myfunc_47_tid_449 <= 0;
      _th_myfunc_47_tid_450 <= 0;
      _th_myfunc_47_time_451 <= 0;
      _th_myfunc_47_i_452 <= 0;
    end else begin
      case(th_myfunc_47)
        th_myfunc_47_init: begin
          if(_th_myfunc_start[47] && (th_blink == 10)) begin
            _th_myfunc_47_called <= 1;
          end 
          if(_th_myfunc_start[47] && (th_blink == 10)) begin
            _th_myfunc_47_tid_449 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[47]) begin
            th_myfunc_47 <= th_myfunc_47_1;
          end 
        end
        th_myfunc_47_1: begin
          _th_myfunc_47_tid_450 <= _th_myfunc_47_tid_449;
          th_myfunc_47 <= th_myfunc_47_2;
        end
        th_myfunc_47_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 47)) begin
            th_myfunc_47 <= th_myfunc_47_3;
          end 
        end
        th_myfunc_47_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 47))) begin
            th_myfunc_47 <= th_myfunc_47_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 47)) begin
            th_myfunc_47 <= th_myfunc_47_4;
          end 
        end
        th_myfunc_47_4: begin
          $display("Thread %d Lock", _th_myfunc_47_tid_450);
          th_myfunc_47 <= th_myfunc_47_5;
        end
        th_myfunc_47_5: begin
          _th_myfunc_47_time_451 <= sw;
          th_myfunc_47 <= th_myfunc_47_6;
        end
        th_myfunc_47_6: begin
          _th_myfunc_47_i_452 <= 0;
          th_myfunc_47 <= th_myfunc_47_7;
        end
        th_myfunc_47_7: begin
          if(_th_myfunc_47_i_452 < _th_myfunc_47_time_451) begin
            th_myfunc_47 <= th_myfunc_47_8;
          end else begin
            th_myfunc_47 <= th_myfunc_47_9;
          end
        end
        th_myfunc_47_8: begin
          _th_myfunc_47_i_452 <= _th_myfunc_47_i_452 + 1;
          th_myfunc_47 <= th_myfunc_47_7;
        end
        th_myfunc_47_9: begin
          th_myfunc_47 <= th_myfunc_47_10;
        end
        th_myfunc_47_10: begin
          $display("Thread %d count = %d", _th_myfunc_47_tid_450, count);
          th_myfunc_47 <= th_myfunc_47_11;
        end
        th_myfunc_47_11: begin
          th_myfunc_47 <= th_myfunc_47_12;
        end
        th_myfunc_47_12: begin
          $display("Thread %d Unlock", _th_myfunc_47_tid_450);
          th_myfunc_47 <= th_myfunc_47_13;
        end
        th_myfunc_47_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 47)) begin
            _th_myfunc_47_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 47)) begin
            th_myfunc_47 <= th_myfunc_47_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_48_1 = 1;
  localparam th_myfunc_48_2 = 2;
  localparam th_myfunc_48_3 = 3;
  localparam th_myfunc_48_4 = 4;
  localparam th_myfunc_48_5 = 5;
  localparam th_myfunc_48_6 = 6;
  localparam th_myfunc_48_7 = 7;
  localparam th_myfunc_48_8 = 8;
  localparam th_myfunc_48_9 = 9;
  localparam th_myfunc_48_10 = 10;
  localparam th_myfunc_48_11 = 11;
  localparam th_myfunc_48_12 = 12;
  localparam th_myfunc_48_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_48 <= th_myfunc_48_init;
      _th_myfunc_48_called <= 0;
      _th_myfunc_48_tid_453 <= 0;
      _th_myfunc_48_tid_454 <= 0;
      _th_myfunc_48_time_455 <= 0;
      _th_myfunc_48_i_456 <= 0;
    end else begin
      case(th_myfunc_48)
        th_myfunc_48_init: begin
          if(_th_myfunc_start[48] && (th_blink == 10)) begin
            _th_myfunc_48_called <= 1;
          end 
          if(_th_myfunc_start[48] && (th_blink == 10)) begin
            _th_myfunc_48_tid_453 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[48]) begin
            th_myfunc_48 <= th_myfunc_48_1;
          end 
        end
        th_myfunc_48_1: begin
          _th_myfunc_48_tid_454 <= _th_myfunc_48_tid_453;
          th_myfunc_48 <= th_myfunc_48_2;
        end
        th_myfunc_48_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 48)) begin
            th_myfunc_48 <= th_myfunc_48_3;
          end 
        end
        th_myfunc_48_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 48))) begin
            th_myfunc_48 <= th_myfunc_48_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 48)) begin
            th_myfunc_48 <= th_myfunc_48_4;
          end 
        end
        th_myfunc_48_4: begin
          $display("Thread %d Lock", _th_myfunc_48_tid_454);
          th_myfunc_48 <= th_myfunc_48_5;
        end
        th_myfunc_48_5: begin
          _th_myfunc_48_time_455 <= sw;
          th_myfunc_48 <= th_myfunc_48_6;
        end
        th_myfunc_48_6: begin
          _th_myfunc_48_i_456 <= 0;
          th_myfunc_48 <= th_myfunc_48_7;
        end
        th_myfunc_48_7: begin
          if(_th_myfunc_48_i_456 < _th_myfunc_48_time_455) begin
            th_myfunc_48 <= th_myfunc_48_8;
          end else begin
            th_myfunc_48 <= th_myfunc_48_9;
          end
        end
        th_myfunc_48_8: begin
          _th_myfunc_48_i_456 <= _th_myfunc_48_i_456 + 1;
          th_myfunc_48 <= th_myfunc_48_7;
        end
        th_myfunc_48_9: begin
          th_myfunc_48 <= th_myfunc_48_10;
        end
        th_myfunc_48_10: begin
          $display("Thread %d count = %d", _th_myfunc_48_tid_454, count);
          th_myfunc_48 <= th_myfunc_48_11;
        end
        th_myfunc_48_11: begin
          th_myfunc_48 <= th_myfunc_48_12;
        end
        th_myfunc_48_12: begin
          $display("Thread %d Unlock", _th_myfunc_48_tid_454);
          th_myfunc_48 <= th_myfunc_48_13;
        end
        th_myfunc_48_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 48)) begin
            _th_myfunc_48_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 48)) begin
            th_myfunc_48 <= th_myfunc_48_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_49_1 = 1;
  localparam th_myfunc_49_2 = 2;
  localparam th_myfunc_49_3 = 3;
  localparam th_myfunc_49_4 = 4;
  localparam th_myfunc_49_5 = 5;
  localparam th_myfunc_49_6 = 6;
  localparam th_myfunc_49_7 = 7;
  localparam th_myfunc_49_8 = 8;
  localparam th_myfunc_49_9 = 9;
  localparam th_myfunc_49_10 = 10;
  localparam th_myfunc_49_11 = 11;
  localparam th_myfunc_49_12 = 12;
  localparam th_myfunc_49_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_49 <= th_myfunc_49_init;
      _th_myfunc_49_called <= 0;
      _th_myfunc_49_tid_457 <= 0;
      _th_myfunc_49_tid_458 <= 0;
      _th_myfunc_49_time_459 <= 0;
      _th_myfunc_49_i_460 <= 0;
    end else begin
      case(th_myfunc_49)
        th_myfunc_49_init: begin
          if(_th_myfunc_start[49] && (th_blink == 10)) begin
            _th_myfunc_49_called <= 1;
          end 
          if(_th_myfunc_start[49] && (th_blink == 10)) begin
            _th_myfunc_49_tid_457 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[49]) begin
            th_myfunc_49 <= th_myfunc_49_1;
          end 
        end
        th_myfunc_49_1: begin
          _th_myfunc_49_tid_458 <= _th_myfunc_49_tid_457;
          th_myfunc_49 <= th_myfunc_49_2;
        end
        th_myfunc_49_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 49)) begin
            th_myfunc_49 <= th_myfunc_49_3;
          end 
        end
        th_myfunc_49_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 49))) begin
            th_myfunc_49 <= th_myfunc_49_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 49)) begin
            th_myfunc_49 <= th_myfunc_49_4;
          end 
        end
        th_myfunc_49_4: begin
          $display("Thread %d Lock", _th_myfunc_49_tid_458);
          th_myfunc_49 <= th_myfunc_49_5;
        end
        th_myfunc_49_5: begin
          _th_myfunc_49_time_459 <= sw;
          th_myfunc_49 <= th_myfunc_49_6;
        end
        th_myfunc_49_6: begin
          _th_myfunc_49_i_460 <= 0;
          th_myfunc_49 <= th_myfunc_49_7;
        end
        th_myfunc_49_7: begin
          if(_th_myfunc_49_i_460 < _th_myfunc_49_time_459) begin
            th_myfunc_49 <= th_myfunc_49_8;
          end else begin
            th_myfunc_49 <= th_myfunc_49_9;
          end
        end
        th_myfunc_49_8: begin
          _th_myfunc_49_i_460 <= _th_myfunc_49_i_460 + 1;
          th_myfunc_49 <= th_myfunc_49_7;
        end
        th_myfunc_49_9: begin
          th_myfunc_49 <= th_myfunc_49_10;
        end
        th_myfunc_49_10: begin
          $display("Thread %d count = %d", _th_myfunc_49_tid_458, count);
          th_myfunc_49 <= th_myfunc_49_11;
        end
        th_myfunc_49_11: begin
          th_myfunc_49 <= th_myfunc_49_12;
        end
        th_myfunc_49_12: begin
          $display("Thread %d Unlock", _th_myfunc_49_tid_458);
          th_myfunc_49 <= th_myfunc_49_13;
        end
        th_myfunc_49_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 49)) begin
            _th_myfunc_49_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 49)) begin
            th_myfunc_49 <= th_myfunc_49_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_50_1 = 1;
  localparam th_myfunc_50_2 = 2;
  localparam th_myfunc_50_3 = 3;
  localparam th_myfunc_50_4 = 4;
  localparam th_myfunc_50_5 = 5;
  localparam th_myfunc_50_6 = 6;
  localparam th_myfunc_50_7 = 7;
  localparam th_myfunc_50_8 = 8;
  localparam th_myfunc_50_9 = 9;
  localparam th_myfunc_50_10 = 10;
  localparam th_myfunc_50_11 = 11;
  localparam th_myfunc_50_12 = 12;
  localparam th_myfunc_50_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_50 <= th_myfunc_50_init;
      _th_myfunc_50_called <= 0;
      _th_myfunc_50_tid_461 <= 0;
      _th_myfunc_50_tid_462 <= 0;
      _th_myfunc_50_time_463 <= 0;
      _th_myfunc_50_i_464 <= 0;
    end else begin
      case(th_myfunc_50)
        th_myfunc_50_init: begin
          if(_th_myfunc_start[50] && (th_blink == 10)) begin
            _th_myfunc_50_called <= 1;
          end 
          if(_th_myfunc_start[50] && (th_blink == 10)) begin
            _th_myfunc_50_tid_461 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[50]) begin
            th_myfunc_50 <= th_myfunc_50_1;
          end 
        end
        th_myfunc_50_1: begin
          _th_myfunc_50_tid_462 <= _th_myfunc_50_tid_461;
          th_myfunc_50 <= th_myfunc_50_2;
        end
        th_myfunc_50_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 50)) begin
            th_myfunc_50 <= th_myfunc_50_3;
          end 
        end
        th_myfunc_50_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 50))) begin
            th_myfunc_50 <= th_myfunc_50_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 50)) begin
            th_myfunc_50 <= th_myfunc_50_4;
          end 
        end
        th_myfunc_50_4: begin
          $display("Thread %d Lock", _th_myfunc_50_tid_462);
          th_myfunc_50 <= th_myfunc_50_5;
        end
        th_myfunc_50_5: begin
          _th_myfunc_50_time_463 <= sw;
          th_myfunc_50 <= th_myfunc_50_6;
        end
        th_myfunc_50_6: begin
          _th_myfunc_50_i_464 <= 0;
          th_myfunc_50 <= th_myfunc_50_7;
        end
        th_myfunc_50_7: begin
          if(_th_myfunc_50_i_464 < _th_myfunc_50_time_463) begin
            th_myfunc_50 <= th_myfunc_50_8;
          end else begin
            th_myfunc_50 <= th_myfunc_50_9;
          end
        end
        th_myfunc_50_8: begin
          _th_myfunc_50_i_464 <= _th_myfunc_50_i_464 + 1;
          th_myfunc_50 <= th_myfunc_50_7;
        end
        th_myfunc_50_9: begin
          th_myfunc_50 <= th_myfunc_50_10;
        end
        th_myfunc_50_10: begin
          $display("Thread %d count = %d", _th_myfunc_50_tid_462, count);
          th_myfunc_50 <= th_myfunc_50_11;
        end
        th_myfunc_50_11: begin
          th_myfunc_50 <= th_myfunc_50_12;
        end
        th_myfunc_50_12: begin
          $display("Thread %d Unlock", _th_myfunc_50_tid_462);
          th_myfunc_50 <= th_myfunc_50_13;
        end
        th_myfunc_50_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 50)) begin
            _th_myfunc_50_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 50)) begin
            th_myfunc_50 <= th_myfunc_50_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_51_1 = 1;
  localparam th_myfunc_51_2 = 2;
  localparam th_myfunc_51_3 = 3;
  localparam th_myfunc_51_4 = 4;
  localparam th_myfunc_51_5 = 5;
  localparam th_myfunc_51_6 = 6;
  localparam th_myfunc_51_7 = 7;
  localparam th_myfunc_51_8 = 8;
  localparam th_myfunc_51_9 = 9;
  localparam th_myfunc_51_10 = 10;
  localparam th_myfunc_51_11 = 11;
  localparam th_myfunc_51_12 = 12;
  localparam th_myfunc_51_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_51 <= th_myfunc_51_init;
      _th_myfunc_51_called <= 0;
      _th_myfunc_51_tid_465 <= 0;
      _th_myfunc_51_tid_466 <= 0;
      _th_myfunc_51_time_467 <= 0;
      _th_myfunc_51_i_468 <= 0;
    end else begin
      case(th_myfunc_51)
        th_myfunc_51_init: begin
          if(_th_myfunc_start[51] && (th_blink == 10)) begin
            _th_myfunc_51_called <= 1;
          end 
          if(_th_myfunc_start[51] && (th_blink == 10)) begin
            _th_myfunc_51_tid_465 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[51]) begin
            th_myfunc_51 <= th_myfunc_51_1;
          end 
        end
        th_myfunc_51_1: begin
          _th_myfunc_51_tid_466 <= _th_myfunc_51_tid_465;
          th_myfunc_51 <= th_myfunc_51_2;
        end
        th_myfunc_51_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 51)) begin
            th_myfunc_51 <= th_myfunc_51_3;
          end 
        end
        th_myfunc_51_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 51))) begin
            th_myfunc_51 <= th_myfunc_51_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 51)) begin
            th_myfunc_51 <= th_myfunc_51_4;
          end 
        end
        th_myfunc_51_4: begin
          $display("Thread %d Lock", _th_myfunc_51_tid_466);
          th_myfunc_51 <= th_myfunc_51_5;
        end
        th_myfunc_51_5: begin
          _th_myfunc_51_time_467 <= sw;
          th_myfunc_51 <= th_myfunc_51_6;
        end
        th_myfunc_51_6: begin
          _th_myfunc_51_i_468 <= 0;
          th_myfunc_51 <= th_myfunc_51_7;
        end
        th_myfunc_51_7: begin
          if(_th_myfunc_51_i_468 < _th_myfunc_51_time_467) begin
            th_myfunc_51 <= th_myfunc_51_8;
          end else begin
            th_myfunc_51 <= th_myfunc_51_9;
          end
        end
        th_myfunc_51_8: begin
          _th_myfunc_51_i_468 <= _th_myfunc_51_i_468 + 1;
          th_myfunc_51 <= th_myfunc_51_7;
        end
        th_myfunc_51_9: begin
          th_myfunc_51 <= th_myfunc_51_10;
        end
        th_myfunc_51_10: begin
          $display("Thread %d count = %d", _th_myfunc_51_tid_466, count);
          th_myfunc_51 <= th_myfunc_51_11;
        end
        th_myfunc_51_11: begin
          th_myfunc_51 <= th_myfunc_51_12;
        end
        th_myfunc_51_12: begin
          $display("Thread %d Unlock", _th_myfunc_51_tid_466);
          th_myfunc_51 <= th_myfunc_51_13;
        end
        th_myfunc_51_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 51)) begin
            _th_myfunc_51_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 51)) begin
            th_myfunc_51 <= th_myfunc_51_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_52_1 = 1;
  localparam th_myfunc_52_2 = 2;
  localparam th_myfunc_52_3 = 3;
  localparam th_myfunc_52_4 = 4;
  localparam th_myfunc_52_5 = 5;
  localparam th_myfunc_52_6 = 6;
  localparam th_myfunc_52_7 = 7;
  localparam th_myfunc_52_8 = 8;
  localparam th_myfunc_52_9 = 9;
  localparam th_myfunc_52_10 = 10;
  localparam th_myfunc_52_11 = 11;
  localparam th_myfunc_52_12 = 12;
  localparam th_myfunc_52_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_52 <= th_myfunc_52_init;
      _th_myfunc_52_called <= 0;
      _th_myfunc_52_tid_469 <= 0;
      _th_myfunc_52_tid_470 <= 0;
      _th_myfunc_52_time_471 <= 0;
      _th_myfunc_52_i_472 <= 0;
    end else begin
      case(th_myfunc_52)
        th_myfunc_52_init: begin
          if(_th_myfunc_start[52] && (th_blink == 10)) begin
            _th_myfunc_52_called <= 1;
          end 
          if(_th_myfunc_start[52] && (th_blink == 10)) begin
            _th_myfunc_52_tid_469 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[52]) begin
            th_myfunc_52 <= th_myfunc_52_1;
          end 
        end
        th_myfunc_52_1: begin
          _th_myfunc_52_tid_470 <= _th_myfunc_52_tid_469;
          th_myfunc_52 <= th_myfunc_52_2;
        end
        th_myfunc_52_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 52)) begin
            th_myfunc_52 <= th_myfunc_52_3;
          end 
        end
        th_myfunc_52_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 52))) begin
            th_myfunc_52 <= th_myfunc_52_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 52)) begin
            th_myfunc_52 <= th_myfunc_52_4;
          end 
        end
        th_myfunc_52_4: begin
          $display("Thread %d Lock", _th_myfunc_52_tid_470);
          th_myfunc_52 <= th_myfunc_52_5;
        end
        th_myfunc_52_5: begin
          _th_myfunc_52_time_471 <= sw;
          th_myfunc_52 <= th_myfunc_52_6;
        end
        th_myfunc_52_6: begin
          _th_myfunc_52_i_472 <= 0;
          th_myfunc_52 <= th_myfunc_52_7;
        end
        th_myfunc_52_7: begin
          if(_th_myfunc_52_i_472 < _th_myfunc_52_time_471) begin
            th_myfunc_52 <= th_myfunc_52_8;
          end else begin
            th_myfunc_52 <= th_myfunc_52_9;
          end
        end
        th_myfunc_52_8: begin
          _th_myfunc_52_i_472 <= _th_myfunc_52_i_472 + 1;
          th_myfunc_52 <= th_myfunc_52_7;
        end
        th_myfunc_52_9: begin
          th_myfunc_52 <= th_myfunc_52_10;
        end
        th_myfunc_52_10: begin
          $display("Thread %d count = %d", _th_myfunc_52_tid_470, count);
          th_myfunc_52 <= th_myfunc_52_11;
        end
        th_myfunc_52_11: begin
          th_myfunc_52 <= th_myfunc_52_12;
        end
        th_myfunc_52_12: begin
          $display("Thread %d Unlock", _th_myfunc_52_tid_470);
          th_myfunc_52 <= th_myfunc_52_13;
        end
        th_myfunc_52_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 52)) begin
            _th_myfunc_52_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 52)) begin
            th_myfunc_52 <= th_myfunc_52_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_53_1 = 1;
  localparam th_myfunc_53_2 = 2;
  localparam th_myfunc_53_3 = 3;
  localparam th_myfunc_53_4 = 4;
  localparam th_myfunc_53_5 = 5;
  localparam th_myfunc_53_6 = 6;
  localparam th_myfunc_53_7 = 7;
  localparam th_myfunc_53_8 = 8;
  localparam th_myfunc_53_9 = 9;
  localparam th_myfunc_53_10 = 10;
  localparam th_myfunc_53_11 = 11;
  localparam th_myfunc_53_12 = 12;
  localparam th_myfunc_53_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_53 <= th_myfunc_53_init;
      _th_myfunc_53_called <= 0;
      _th_myfunc_53_tid_473 <= 0;
      _th_myfunc_53_tid_474 <= 0;
      _th_myfunc_53_time_475 <= 0;
      _th_myfunc_53_i_476 <= 0;
    end else begin
      case(th_myfunc_53)
        th_myfunc_53_init: begin
          if(_th_myfunc_start[53] && (th_blink == 10)) begin
            _th_myfunc_53_called <= 1;
          end 
          if(_th_myfunc_start[53] && (th_blink == 10)) begin
            _th_myfunc_53_tid_473 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[53]) begin
            th_myfunc_53 <= th_myfunc_53_1;
          end 
        end
        th_myfunc_53_1: begin
          _th_myfunc_53_tid_474 <= _th_myfunc_53_tid_473;
          th_myfunc_53 <= th_myfunc_53_2;
        end
        th_myfunc_53_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 53)) begin
            th_myfunc_53 <= th_myfunc_53_3;
          end 
        end
        th_myfunc_53_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 53))) begin
            th_myfunc_53 <= th_myfunc_53_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 53)) begin
            th_myfunc_53 <= th_myfunc_53_4;
          end 
        end
        th_myfunc_53_4: begin
          $display("Thread %d Lock", _th_myfunc_53_tid_474);
          th_myfunc_53 <= th_myfunc_53_5;
        end
        th_myfunc_53_5: begin
          _th_myfunc_53_time_475 <= sw;
          th_myfunc_53 <= th_myfunc_53_6;
        end
        th_myfunc_53_6: begin
          _th_myfunc_53_i_476 <= 0;
          th_myfunc_53 <= th_myfunc_53_7;
        end
        th_myfunc_53_7: begin
          if(_th_myfunc_53_i_476 < _th_myfunc_53_time_475) begin
            th_myfunc_53 <= th_myfunc_53_8;
          end else begin
            th_myfunc_53 <= th_myfunc_53_9;
          end
        end
        th_myfunc_53_8: begin
          _th_myfunc_53_i_476 <= _th_myfunc_53_i_476 + 1;
          th_myfunc_53 <= th_myfunc_53_7;
        end
        th_myfunc_53_9: begin
          th_myfunc_53 <= th_myfunc_53_10;
        end
        th_myfunc_53_10: begin
          $display("Thread %d count = %d", _th_myfunc_53_tid_474, count);
          th_myfunc_53 <= th_myfunc_53_11;
        end
        th_myfunc_53_11: begin
          th_myfunc_53 <= th_myfunc_53_12;
        end
        th_myfunc_53_12: begin
          $display("Thread %d Unlock", _th_myfunc_53_tid_474);
          th_myfunc_53 <= th_myfunc_53_13;
        end
        th_myfunc_53_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 53)) begin
            _th_myfunc_53_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 53)) begin
            th_myfunc_53 <= th_myfunc_53_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_54_1 = 1;
  localparam th_myfunc_54_2 = 2;
  localparam th_myfunc_54_3 = 3;
  localparam th_myfunc_54_4 = 4;
  localparam th_myfunc_54_5 = 5;
  localparam th_myfunc_54_6 = 6;
  localparam th_myfunc_54_7 = 7;
  localparam th_myfunc_54_8 = 8;
  localparam th_myfunc_54_9 = 9;
  localparam th_myfunc_54_10 = 10;
  localparam th_myfunc_54_11 = 11;
  localparam th_myfunc_54_12 = 12;
  localparam th_myfunc_54_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_54 <= th_myfunc_54_init;
      _th_myfunc_54_called <= 0;
      _th_myfunc_54_tid_477 <= 0;
      _th_myfunc_54_tid_478 <= 0;
      _th_myfunc_54_time_479 <= 0;
      _th_myfunc_54_i_480 <= 0;
    end else begin
      case(th_myfunc_54)
        th_myfunc_54_init: begin
          if(_th_myfunc_start[54] && (th_blink == 10)) begin
            _th_myfunc_54_called <= 1;
          end 
          if(_th_myfunc_start[54] && (th_blink == 10)) begin
            _th_myfunc_54_tid_477 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[54]) begin
            th_myfunc_54 <= th_myfunc_54_1;
          end 
        end
        th_myfunc_54_1: begin
          _th_myfunc_54_tid_478 <= _th_myfunc_54_tid_477;
          th_myfunc_54 <= th_myfunc_54_2;
        end
        th_myfunc_54_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 54)) begin
            th_myfunc_54 <= th_myfunc_54_3;
          end 
        end
        th_myfunc_54_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 54))) begin
            th_myfunc_54 <= th_myfunc_54_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 54)) begin
            th_myfunc_54 <= th_myfunc_54_4;
          end 
        end
        th_myfunc_54_4: begin
          $display("Thread %d Lock", _th_myfunc_54_tid_478);
          th_myfunc_54 <= th_myfunc_54_5;
        end
        th_myfunc_54_5: begin
          _th_myfunc_54_time_479 <= sw;
          th_myfunc_54 <= th_myfunc_54_6;
        end
        th_myfunc_54_6: begin
          _th_myfunc_54_i_480 <= 0;
          th_myfunc_54 <= th_myfunc_54_7;
        end
        th_myfunc_54_7: begin
          if(_th_myfunc_54_i_480 < _th_myfunc_54_time_479) begin
            th_myfunc_54 <= th_myfunc_54_8;
          end else begin
            th_myfunc_54 <= th_myfunc_54_9;
          end
        end
        th_myfunc_54_8: begin
          _th_myfunc_54_i_480 <= _th_myfunc_54_i_480 + 1;
          th_myfunc_54 <= th_myfunc_54_7;
        end
        th_myfunc_54_9: begin
          th_myfunc_54 <= th_myfunc_54_10;
        end
        th_myfunc_54_10: begin
          $display("Thread %d count = %d", _th_myfunc_54_tid_478, count);
          th_myfunc_54 <= th_myfunc_54_11;
        end
        th_myfunc_54_11: begin
          th_myfunc_54 <= th_myfunc_54_12;
        end
        th_myfunc_54_12: begin
          $display("Thread %d Unlock", _th_myfunc_54_tid_478);
          th_myfunc_54 <= th_myfunc_54_13;
        end
        th_myfunc_54_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 54)) begin
            _th_myfunc_54_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 54)) begin
            th_myfunc_54 <= th_myfunc_54_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_55_1 = 1;
  localparam th_myfunc_55_2 = 2;
  localparam th_myfunc_55_3 = 3;
  localparam th_myfunc_55_4 = 4;
  localparam th_myfunc_55_5 = 5;
  localparam th_myfunc_55_6 = 6;
  localparam th_myfunc_55_7 = 7;
  localparam th_myfunc_55_8 = 8;
  localparam th_myfunc_55_9 = 9;
  localparam th_myfunc_55_10 = 10;
  localparam th_myfunc_55_11 = 11;
  localparam th_myfunc_55_12 = 12;
  localparam th_myfunc_55_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_55 <= th_myfunc_55_init;
      _th_myfunc_55_called <= 0;
      _th_myfunc_55_tid_481 <= 0;
      _th_myfunc_55_tid_482 <= 0;
      _th_myfunc_55_time_483 <= 0;
      _th_myfunc_55_i_484 <= 0;
    end else begin
      case(th_myfunc_55)
        th_myfunc_55_init: begin
          if(_th_myfunc_start[55] && (th_blink == 10)) begin
            _th_myfunc_55_called <= 1;
          end 
          if(_th_myfunc_start[55] && (th_blink == 10)) begin
            _th_myfunc_55_tid_481 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[55]) begin
            th_myfunc_55 <= th_myfunc_55_1;
          end 
        end
        th_myfunc_55_1: begin
          _th_myfunc_55_tid_482 <= _th_myfunc_55_tid_481;
          th_myfunc_55 <= th_myfunc_55_2;
        end
        th_myfunc_55_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 55)) begin
            th_myfunc_55 <= th_myfunc_55_3;
          end 
        end
        th_myfunc_55_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 55))) begin
            th_myfunc_55 <= th_myfunc_55_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 55)) begin
            th_myfunc_55 <= th_myfunc_55_4;
          end 
        end
        th_myfunc_55_4: begin
          $display("Thread %d Lock", _th_myfunc_55_tid_482);
          th_myfunc_55 <= th_myfunc_55_5;
        end
        th_myfunc_55_5: begin
          _th_myfunc_55_time_483 <= sw;
          th_myfunc_55 <= th_myfunc_55_6;
        end
        th_myfunc_55_6: begin
          _th_myfunc_55_i_484 <= 0;
          th_myfunc_55 <= th_myfunc_55_7;
        end
        th_myfunc_55_7: begin
          if(_th_myfunc_55_i_484 < _th_myfunc_55_time_483) begin
            th_myfunc_55 <= th_myfunc_55_8;
          end else begin
            th_myfunc_55 <= th_myfunc_55_9;
          end
        end
        th_myfunc_55_8: begin
          _th_myfunc_55_i_484 <= _th_myfunc_55_i_484 + 1;
          th_myfunc_55 <= th_myfunc_55_7;
        end
        th_myfunc_55_9: begin
          th_myfunc_55 <= th_myfunc_55_10;
        end
        th_myfunc_55_10: begin
          $display("Thread %d count = %d", _th_myfunc_55_tid_482, count);
          th_myfunc_55 <= th_myfunc_55_11;
        end
        th_myfunc_55_11: begin
          th_myfunc_55 <= th_myfunc_55_12;
        end
        th_myfunc_55_12: begin
          $display("Thread %d Unlock", _th_myfunc_55_tid_482);
          th_myfunc_55 <= th_myfunc_55_13;
        end
        th_myfunc_55_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 55)) begin
            _th_myfunc_55_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 55)) begin
            th_myfunc_55 <= th_myfunc_55_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_56_1 = 1;
  localparam th_myfunc_56_2 = 2;
  localparam th_myfunc_56_3 = 3;
  localparam th_myfunc_56_4 = 4;
  localparam th_myfunc_56_5 = 5;
  localparam th_myfunc_56_6 = 6;
  localparam th_myfunc_56_7 = 7;
  localparam th_myfunc_56_8 = 8;
  localparam th_myfunc_56_9 = 9;
  localparam th_myfunc_56_10 = 10;
  localparam th_myfunc_56_11 = 11;
  localparam th_myfunc_56_12 = 12;
  localparam th_myfunc_56_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_56 <= th_myfunc_56_init;
      _th_myfunc_56_called <= 0;
      _th_myfunc_56_tid_485 <= 0;
      _th_myfunc_56_tid_486 <= 0;
      _th_myfunc_56_time_487 <= 0;
      _th_myfunc_56_i_488 <= 0;
    end else begin
      case(th_myfunc_56)
        th_myfunc_56_init: begin
          if(_th_myfunc_start[56] && (th_blink == 10)) begin
            _th_myfunc_56_called <= 1;
          end 
          if(_th_myfunc_start[56] && (th_blink == 10)) begin
            _th_myfunc_56_tid_485 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[56]) begin
            th_myfunc_56 <= th_myfunc_56_1;
          end 
        end
        th_myfunc_56_1: begin
          _th_myfunc_56_tid_486 <= _th_myfunc_56_tid_485;
          th_myfunc_56 <= th_myfunc_56_2;
        end
        th_myfunc_56_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 56)) begin
            th_myfunc_56 <= th_myfunc_56_3;
          end 
        end
        th_myfunc_56_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 56))) begin
            th_myfunc_56 <= th_myfunc_56_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 56)) begin
            th_myfunc_56 <= th_myfunc_56_4;
          end 
        end
        th_myfunc_56_4: begin
          $display("Thread %d Lock", _th_myfunc_56_tid_486);
          th_myfunc_56 <= th_myfunc_56_5;
        end
        th_myfunc_56_5: begin
          _th_myfunc_56_time_487 <= sw;
          th_myfunc_56 <= th_myfunc_56_6;
        end
        th_myfunc_56_6: begin
          _th_myfunc_56_i_488 <= 0;
          th_myfunc_56 <= th_myfunc_56_7;
        end
        th_myfunc_56_7: begin
          if(_th_myfunc_56_i_488 < _th_myfunc_56_time_487) begin
            th_myfunc_56 <= th_myfunc_56_8;
          end else begin
            th_myfunc_56 <= th_myfunc_56_9;
          end
        end
        th_myfunc_56_8: begin
          _th_myfunc_56_i_488 <= _th_myfunc_56_i_488 + 1;
          th_myfunc_56 <= th_myfunc_56_7;
        end
        th_myfunc_56_9: begin
          th_myfunc_56 <= th_myfunc_56_10;
        end
        th_myfunc_56_10: begin
          $display("Thread %d count = %d", _th_myfunc_56_tid_486, count);
          th_myfunc_56 <= th_myfunc_56_11;
        end
        th_myfunc_56_11: begin
          th_myfunc_56 <= th_myfunc_56_12;
        end
        th_myfunc_56_12: begin
          $display("Thread %d Unlock", _th_myfunc_56_tid_486);
          th_myfunc_56 <= th_myfunc_56_13;
        end
        th_myfunc_56_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 56)) begin
            _th_myfunc_56_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 56)) begin
            th_myfunc_56 <= th_myfunc_56_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_57_1 = 1;
  localparam th_myfunc_57_2 = 2;
  localparam th_myfunc_57_3 = 3;
  localparam th_myfunc_57_4 = 4;
  localparam th_myfunc_57_5 = 5;
  localparam th_myfunc_57_6 = 6;
  localparam th_myfunc_57_7 = 7;
  localparam th_myfunc_57_8 = 8;
  localparam th_myfunc_57_9 = 9;
  localparam th_myfunc_57_10 = 10;
  localparam th_myfunc_57_11 = 11;
  localparam th_myfunc_57_12 = 12;
  localparam th_myfunc_57_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_57 <= th_myfunc_57_init;
      _th_myfunc_57_called <= 0;
      _th_myfunc_57_tid_489 <= 0;
      _th_myfunc_57_tid_490 <= 0;
      _th_myfunc_57_time_491 <= 0;
      _th_myfunc_57_i_492 <= 0;
    end else begin
      case(th_myfunc_57)
        th_myfunc_57_init: begin
          if(_th_myfunc_start[57] && (th_blink == 10)) begin
            _th_myfunc_57_called <= 1;
          end 
          if(_th_myfunc_start[57] && (th_blink == 10)) begin
            _th_myfunc_57_tid_489 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[57]) begin
            th_myfunc_57 <= th_myfunc_57_1;
          end 
        end
        th_myfunc_57_1: begin
          _th_myfunc_57_tid_490 <= _th_myfunc_57_tid_489;
          th_myfunc_57 <= th_myfunc_57_2;
        end
        th_myfunc_57_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 57)) begin
            th_myfunc_57 <= th_myfunc_57_3;
          end 
        end
        th_myfunc_57_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 57))) begin
            th_myfunc_57 <= th_myfunc_57_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 57)) begin
            th_myfunc_57 <= th_myfunc_57_4;
          end 
        end
        th_myfunc_57_4: begin
          $display("Thread %d Lock", _th_myfunc_57_tid_490);
          th_myfunc_57 <= th_myfunc_57_5;
        end
        th_myfunc_57_5: begin
          _th_myfunc_57_time_491 <= sw;
          th_myfunc_57 <= th_myfunc_57_6;
        end
        th_myfunc_57_6: begin
          _th_myfunc_57_i_492 <= 0;
          th_myfunc_57 <= th_myfunc_57_7;
        end
        th_myfunc_57_7: begin
          if(_th_myfunc_57_i_492 < _th_myfunc_57_time_491) begin
            th_myfunc_57 <= th_myfunc_57_8;
          end else begin
            th_myfunc_57 <= th_myfunc_57_9;
          end
        end
        th_myfunc_57_8: begin
          _th_myfunc_57_i_492 <= _th_myfunc_57_i_492 + 1;
          th_myfunc_57 <= th_myfunc_57_7;
        end
        th_myfunc_57_9: begin
          th_myfunc_57 <= th_myfunc_57_10;
        end
        th_myfunc_57_10: begin
          $display("Thread %d count = %d", _th_myfunc_57_tid_490, count);
          th_myfunc_57 <= th_myfunc_57_11;
        end
        th_myfunc_57_11: begin
          th_myfunc_57 <= th_myfunc_57_12;
        end
        th_myfunc_57_12: begin
          $display("Thread %d Unlock", _th_myfunc_57_tid_490);
          th_myfunc_57 <= th_myfunc_57_13;
        end
        th_myfunc_57_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 57)) begin
            _th_myfunc_57_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 57)) begin
            th_myfunc_57 <= th_myfunc_57_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_58_1 = 1;
  localparam th_myfunc_58_2 = 2;
  localparam th_myfunc_58_3 = 3;
  localparam th_myfunc_58_4 = 4;
  localparam th_myfunc_58_5 = 5;
  localparam th_myfunc_58_6 = 6;
  localparam th_myfunc_58_7 = 7;
  localparam th_myfunc_58_8 = 8;
  localparam th_myfunc_58_9 = 9;
  localparam th_myfunc_58_10 = 10;
  localparam th_myfunc_58_11 = 11;
  localparam th_myfunc_58_12 = 12;
  localparam th_myfunc_58_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_58 <= th_myfunc_58_init;
      _th_myfunc_58_called <= 0;
      _th_myfunc_58_tid_493 <= 0;
      _th_myfunc_58_tid_494 <= 0;
      _th_myfunc_58_time_495 <= 0;
      _th_myfunc_58_i_496 <= 0;
    end else begin
      case(th_myfunc_58)
        th_myfunc_58_init: begin
          if(_th_myfunc_start[58] && (th_blink == 10)) begin
            _th_myfunc_58_called <= 1;
          end 
          if(_th_myfunc_start[58] && (th_blink == 10)) begin
            _th_myfunc_58_tid_493 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[58]) begin
            th_myfunc_58 <= th_myfunc_58_1;
          end 
        end
        th_myfunc_58_1: begin
          _th_myfunc_58_tid_494 <= _th_myfunc_58_tid_493;
          th_myfunc_58 <= th_myfunc_58_2;
        end
        th_myfunc_58_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 58)) begin
            th_myfunc_58 <= th_myfunc_58_3;
          end 
        end
        th_myfunc_58_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 58))) begin
            th_myfunc_58 <= th_myfunc_58_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 58)) begin
            th_myfunc_58 <= th_myfunc_58_4;
          end 
        end
        th_myfunc_58_4: begin
          $display("Thread %d Lock", _th_myfunc_58_tid_494);
          th_myfunc_58 <= th_myfunc_58_5;
        end
        th_myfunc_58_5: begin
          _th_myfunc_58_time_495 <= sw;
          th_myfunc_58 <= th_myfunc_58_6;
        end
        th_myfunc_58_6: begin
          _th_myfunc_58_i_496 <= 0;
          th_myfunc_58 <= th_myfunc_58_7;
        end
        th_myfunc_58_7: begin
          if(_th_myfunc_58_i_496 < _th_myfunc_58_time_495) begin
            th_myfunc_58 <= th_myfunc_58_8;
          end else begin
            th_myfunc_58 <= th_myfunc_58_9;
          end
        end
        th_myfunc_58_8: begin
          _th_myfunc_58_i_496 <= _th_myfunc_58_i_496 + 1;
          th_myfunc_58 <= th_myfunc_58_7;
        end
        th_myfunc_58_9: begin
          th_myfunc_58 <= th_myfunc_58_10;
        end
        th_myfunc_58_10: begin
          $display("Thread %d count = %d", _th_myfunc_58_tid_494, count);
          th_myfunc_58 <= th_myfunc_58_11;
        end
        th_myfunc_58_11: begin
          th_myfunc_58 <= th_myfunc_58_12;
        end
        th_myfunc_58_12: begin
          $display("Thread %d Unlock", _th_myfunc_58_tid_494);
          th_myfunc_58 <= th_myfunc_58_13;
        end
        th_myfunc_58_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 58)) begin
            _th_myfunc_58_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 58)) begin
            th_myfunc_58 <= th_myfunc_58_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_59_1 = 1;
  localparam th_myfunc_59_2 = 2;
  localparam th_myfunc_59_3 = 3;
  localparam th_myfunc_59_4 = 4;
  localparam th_myfunc_59_5 = 5;
  localparam th_myfunc_59_6 = 6;
  localparam th_myfunc_59_7 = 7;
  localparam th_myfunc_59_8 = 8;
  localparam th_myfunc_59_9 = 9;
  localparam th_myfunc_59_10 = 10;
  localparam th_myfunc_59_11 = 11;
  localparam th_myfunc_59_12 = 12;
  localparam th_myfunc_59_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_59 <= th_myfunc_59_init;
      _th_myfunc_59_called <= 0;
      _th_myfunc_59_tid_497 <= 0;
      _th_myfunc_59_tid_498 <= 0;
      _th_myfunc_59_time_499 <= 0;
      _th_myfunc_59_i_500 <= 0;
    end else begin
      case(th_myfunc_59)
        th_myfunc_59_init: begin
          if(_th_myfunc_start[59] && (th_blink == 10)) begin
            _th_myfunc_59_called <= 1;
          end 
          if(_th_myfunc_start[59] && (th_blink == 10)) begin
            _th_myfunc_59_tid_497 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[59]) begin
            th_myfunc_59 <= th_myfunc_59_1;
          end 
        end
        th_myfunc_59_1: begin
          _th_myfunc_59_tid_498 <= _th_myfunc_59_tid_497;
          th_myfunc_59 <= th_myfunc_59_2;
        end
        th_myfunc_59_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 59)) begin
            th_myfunc_59 <= th_myfunc_59_3;
          end 
        end
        th_myfunc_59_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 59))) begin
            th_myfunc_59 <= th_myfunc_59_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 59)) begin
            th_myfunc_59 <= th_myfunc_59_4;
          end 
        end
        th_myfunc_59_4: begin
          $display("Thread %d Lock", _th_myfunc_59_tid_498);
          th_myfunc_59 <= th_myfunc_59_5;
        end
        th_myfunc_59_5: begin
          _th_myfunc_59_time_499 <= sw;
          th_myfunc_59 <= th_myfunc_59_6;
        end
        th_myfunc_59_6: begin
          _th_myfunc_59_i_500 <= 0;
          th_myfunc_59 <= th_myfunc_59_7;
        end
        th_myfunc_59_7: begin
          if(_th_myfunc_59_i_500 < _th_myfunc_59_time_499) begin
            th_myfunc_59 <= th_myfunc_59_8;
          end else begin
            th_myfunc_59 <= th_myfunc_59_9;
          end
        end
        th_myfunc_59_8: begin
          _th_myfunc_59_i_500 <= _th_myfunc_59_i_500 + 1;
          th_myfunc_59 <= th_myfunc_59_7;
        end
        th_myfunc_59_9: begin
          th_myfunc_59 <= th_myfunc_59_10;
        end
        th_myfunc_59_10: begin
          $display("Thread %d count = %d", _th_myfunc_59_tid_498, count);
          th_myfunc_59 <= th_myfunc_59_11;
        end
        th_myfunc_59_11: begin
          th_myfunc_59 <= th_myfunc_59_12;
        end
        th_myfunc_59_12: begin
          $display("Thread %d Unlock", _th_myfunc_59_tid_498);
          th_myfunc_59 <= th_myfunc_59_13;
        end
        th_myfunc_59_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 59)) begin
            _th_myfunc_59_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 59)) begin
            th_myfunc_59 <= th_myfunc_59_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_60_1 = 1;
  localparam th_myfunc_60_2 = 2;
  localparam th_myfunc_60_3 = 3;
  localparam th_myfunc_60_4 = 4;
  localparam th_myfunc_60_5 = 5;
  localparam th_myfunc_60_6 = 6;
  localparam th_myfunc_60_7 = 7;
  localparam th_myfunc_60_8 = 8;
  localparam th_myfunc_60_9 = 9;
  localparam th_myfunc_60_10 = 10;
  localparam th_myfunc_60_11 = 11;
  localparam th_myfunc_60_12 = 12;
  localparam th_myfunc_60_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_60 <= th_myfunc_60_init;
      _th_myfunc_60_called <= 0;
      _th_myfunc_60_tid_501 <= 0;
      _th_myfunc_60_tid_502 <= 0;
      _th_myfunc_60_time_503 <= 0;
      _th_myfunc_60_i_504 <= 0;
    end else begin
      case(th_myfunc_60)
        th_myfunc_60_init: begin
          if(_th_myfunc_start[60] && (th_blink == 10)) begin
            _th_myfunc_60_called <= 1;
          end 
          if(_th_myfunc_start[60] && (th_blink == 10)) begin
            _th_myfunc_60_tid_501 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[60]) begin
            th_myfunc_60 <= th_myfunc_60_1;
          end 
        end
        th_myfunc_60_1: begin
          _th_myfunc_60_tid_502 <= _th_myfunc_60_tid_501;
          th_myfunc_60 <= th_myfunc_60_2;
        end
        th_myfunc_60_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 60)) begin
            th_myfunc_60 <= th_myfunc_60_3;
          end 
        end
        th_myfunc_60_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 60))) begin
            th_myfunc_60 <= th_myfunc_60_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 60)) begin
            th_myfunc_60 <= th_myfunc_60_4;
          end 
        end
        th_myfunc_60_4: begin
          $display("Thread %d Lock", _th_myfunc_60_tid_502);
          th_myfunc_60 <= th_myfunc_60_5;
        end
        th_myfunc_60_5: begin
          _th_myfunc_60_time_503 <= sw;
          th_myfunc_60 <= th_myfunc_60_6;
        end
        th_myfunc_60_6: begin
          _th_myfunc_60_i_504 <= 0;
          th_myfunc_60 <= th_myfunc_60_7;
        end
        th_myfunc_60_7: begin
          if(_th_myfunc_60_i_504 < _th_myfunc_60_time_503) begin
            th_myfunc_60 <= th_myfunc_60_8;
          end else begin
            th_myfunc_60 <= th_myfunc_60_9;
          end
        end
        th_myfunc_60_8: begin
          _th_myfunc_60_i_504 <= _th_myfunc_60_i_504 + 1;
          th_myfunc_60 <= th_myfunc_60_7;
        end
        th_myfunc_60_9: begin
          th_myfunc_60 <= th_myfunc_60_10;
        end
        th_myfunc_60_10: begin
          $display("Thread %d count = %d", _th_myfunc_60_tid_502, count);
          th_myfunc_60 <= th_myfunc_60_11;
        end
        th_myfunc_60_11: begin
          th_myfunc_60 <= th_myfunc_60_12;
        end
        th_myfunc_60_12: begin
          $display("Thread %d Unlock", _th_myfunc_60_tid_502);
          th_myfunc_60 <= th_myfunc_60_13;
        end
        th_myfunc_60_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 60)) begin
            _th_myfunc_60_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 60)) begin
            th_myfunc_60 <= th_myfunc_60_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_61_1 = 1;
  localparam th_myfunc_61_2 = 2;
  localparam th_myfunc_61_3 = 3;
  localparam th_myfunc_61_4 = 4;
  localparam th_myfunc_61_5 = 5;
  localparam th_myfunc_61_6 = 6;
  localparam th_myfunc_61_7 = 7;
  localparam th_myfunc_61_8 = 8;
  localparam th_myfunc_61_9 = 9;
  localparam th_myfunc_61_10 = 10;
  localparam th_myfunc_61_11 = 11;
  localparam th_myfunc_61_12 = 12;
  localparam th_myfunc_61_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_61 <= th_myfunc_61_init;
      _th_myfunc_61_called <= 0;
      _th_myfunc_61_tid_505 <= 0;
      _th_myfunc_61_tid_506 <= 0;
      _th_myfunc_61_time_507 <= 0;
      _th_myfunc_61_i_508 <= 0;
    end else begin
      case(th_myfunc_61)
        th_myfunc_61_init: begin
          if(_th_myfunc_start[61] && (th_blink == 10)) begin
            _th_myfunc_61_called <= 1;
          end 
          if(_th_myfunc_start[61] && (th_blink == 10)) begin
            _th_myfunc_61_tid_505 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[61]) begin
            th_myfunc_61 <= th_myfunc_61_1;
          end 
        end
        th_myfunc_61_1: begin
          _th_myfunc_61_tid_506 <= _th_myfunc_61_tid_505;
          th_myfunc_61 <= th_myfunc_61_2;
        end
        th_myfunc_61_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 61)) begin
            th_myfunc_61 <= th_myfunc_61_3;
          end 
        end
        th_myfunc_61_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 61))) begin
            th_myfunc_61 <= th_myfunc_61_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 61)) begin
            th_myfunc_61 <= th_myfunc_61_4;
          end 
        end
        th_myfunc_61_4: begin
          $display("Thread %d Lock", _th_myfunc_61_tid_506);
          th_myfunc_61 <= th_myfunc_61_5;
        end
        th_myfunc_61_5: begin
          _th_myfunc_61_time_507 <= sw;
          th_myfunc_61 <= th_myfunc_61_6;
        end
        th_myfunc_61_6: begin
          _th_myfunc_61_i_508 <= 0;
          th_myfunc_61 <= th_myfunc_61_7;
        end
        th_myfunc_61_7: begin
          if(_th_myfunc_61_i_508 < _th_myfunc_61_time_507) begin
            th_myfunc_61 <= th_myfunc_61_8;
          end else begin
            th_myfunc_61 <= th_myfunc_61_9;
          end
        end
        th_myfunc_61_8: begin
          _th_myfunc_61_i_508 <= _th_myfunc_61_i_508 + 1;
          th_myfunc_61 <= th_myfunc_61_7;
        end
        th_myfunc_61_9: begin
          th_myfunc_61 <= th_myfunc_61_10;
        end
        th_myfunc_61_10: begin
          $display("Thread %d count = %d", _th_myfunc_61_tid_506, count);
          th_myfunc_61 <= th_myfunc_61_11;
        end
        th_myfunc_61_11: begin
          th_myfunc_61 <= th_myfunc_61_12;
        end
        th_myfunc_61_12: begin
          $display("Thread %d Unlock", _th_myfunc_61_tid_506);
          th_myfunc_61 <= th_myfunc_61_13;
        end
        th_myfunc_61_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 61)) begin
            _th_myfunc_61_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 61)) begin
            th_myfunc_61 <= th_myfunc_61_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_62_1 = 1;
  localparam th_myfunc_62_2 = 2;
  localparam th_myfunc_62_3 = 3;
  localparam th_myfunc_62_4 = 4;
  localparam th_myfunc_62_5 = 5;
  localparam th_myfunc_62_6 = 6;
  localparam th_myfunc_62_7 = 7;
  localparam th_myfunc_62_8 = 8;
  localparam th_myfunc_62_9 = 9;
  localparam th_myfunc_62_10 = 10;
  localparam th_myfunc_62_11 = 11;
  localparam th_myfunc_62_12 = 12;
  localparam th_myfunc_62_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_62 <= th_myfunc_62_init;
      _th_myfunc_62_called <= 0;
      _th_myfunc_62_tid_509 <= 0;
      _th_myfunc_62_tid_510 <= 0;
      _th_myfunc_62_time_511 <= 0;
      _th_myfunc_62_i_512 <= 0;
    end else begin
      case(th_myfunc_62)
        th_myfunc_62_init: begin
          if(_th_myfunc_start[62] && (th_blink == 10)) begin
            _th_myfunc_62_called <= 1;
          end 
          if(_th_myfunc_start[62] && (th_blink == 10)) begin
            _th_myfunc_62_tid_509 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[62]) begin
            th_myfunc_62 <= th_myfunc_62_1;
          end 
        end
        th_myfunc_62_1: begin
          _th_myfunc_62_tid_510 <= _th_myfunc_62_tid_509;
          th_myfunc_62 <= th_myfunc_62_2;
        end
        th_myfunc_62_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 62)) begin
            th_myfunc_62 <= th_myfunc_62_3;
          end 
        end
        th_myfunc_62_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 62))) begin
            th_myfunc_62 <= th_myfunc_62_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 62)) begin
            th_myfunc_62 <= th_myfunc_62_4;
          end 
        end
        th_myfunc_62_4: begin
          $display("Thread %d Lock", _th_myfunc_62_tid_510);
          th_myfunc_62 <= th_myfunc_62_5;
        end
        th_myfunc_62_5: begin
          _th_myfunc_62_time_511 <= sw;
          th_myfunc_62 <= th_myfunc_62_6;
        end
        th_myfunc_62_6: begin
          _th_myfunc_62_i_512 <= 0;
          th_myfunc_62 <= th_myfunc_62_7;
        end
        th_myfunc_62_7: begin
          if(_th_myfunc_62_i_512 < _th_myfunc_62_time_511) begin
            th_myfunc_62 <= th_myfunc_62_8;
          end else begin
            th_myfunc_62 <= th_myfunc_62_9;
          end
        end
        th_myfunc_62_8: begin
          _th_myfunc_62_i_512 <= _th_myfunc_62_i_512 + 1;
          th_myfunc_62 <= th_myfunc_62_7;
        end
        th_myfunc_62_9: begin
          th_myfunc_62 <= th_myfunc_62_10;
        end
        th_myfunc_62_10: begin
          $display("Thread %d count = %d", _th_myfunc_62_tid_510, count);
          th_myfunc_62 <= th_myfunc_62_11;
        end
        th_myfunc_62_11: begin
          th_myfunc_62 <= th_myfunc_62_12;
        end
        th_myfunc_62_12: begin
          $display("Thread %d Unlock", _th_myfunc_62_tid_510);
          th_myfunc_62 <= th_myfunc_62_13;
        end
        th_myfunc_62_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 62)) begin
            _th_myfunc_62_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 62)) begin
            th_myfunc_62 <= th_myfunc_62_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_63_1 = 1;
  localparam th_myfunc_63_2 = 2;
  localparam th_myfunc_63_3 = 3;
  localparam th_myfunc_63_4 = 4;
  localparam th_myfunc_63_5 = 5;
  localparam th_myfunc_63_6 = 6;
  localparam th_myfunc_63_7 = 7;
  localparam th_myfunc_63_8 = 8;
  localparam th_myfunc_63_9 = 9;
  localparam th_myfunc_63_10 = 10;
  localparam th_myfunc_63_11 = 11;
  localparam th_myfunc_63_12 = 12;
  localparam th_myfunc_63_13 = 13;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_63 <= th_myfunc_63_init;
      _th_myfunc_63_called <= 0;
      _th_myfunc_63_tid_513 <= 0;
      _th_myfunc_63_tid_514 <= 0;
      _th_myfunc_63_time_515 <= 0;
      _th_myfunc_63_i_516 <= 0;
    end else begin
      case(th_myfunc_63)
        th_myfunc_63_init: begin
          if(_th_myfunc_start[63] && (th_blink == 10)) begin
            _th_myfunc_63_called <= 1;
          end 
          if(_th_myfunc_start[63] && (th_blink == 10)) begin
            _th_myfunc_63_tid_513 <= _th_blink_tid_260;
          end 
          if((th_blink == 10) && _th_myfunc_start[63]) begin
            th_myfunc_63 <= th_myfunc_63_1;
          end 
        end
        th_myfunc_63_1: begin
          _th_myfunc_63_tid_514 <= _th_myfunc_63_tid_513;
          th_myfunc_63 <= th_myfunc_63_2;
        end
        th_myfunc_63_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 63)) begin
            th_myfunc_63 <= th_myfunc_63_3;
          end 
        end
        th_myfunc_63_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 63))) begin
            th_myfunc_63 <= th_myfunc_63_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 63)) begin
            th_myfunc_63 <= th_myfunc_63_4;
          end 
        end
        th_myfunc_63_4: begin
          $display("Thread %d Lock", _th_myfunc_63_tid_514);
          th_myfunc_63 <= th_myfunc_63_5;
        end
        th_myfunc_63_5: begin
          _th_myfunc_63_time_515 <= sw;
          th_myfunc_63 <= th_myfunc_63_6;
        end
        th_myfunc_63_6: begin
          _th_myfunc_63_i_516 <= 0;
          th_myfunc_63 <= th_myfunc_63_7;
        end
        th_myfunc_63_7: begin
          if(_th_myfunc_63_i_516 < _th_myfunc_63_time_515) begin
            th_myfunc_63 <= th_myfunc_63_8;
          end else begin
            th_myfunc_63 <= th_myfunc_63_9;
          end
        end
        th_myfunc_63_8: begin
          _th_myfunc_63_i_516 <= _th_myfunc_63_i_516 + 1;
          th_myfunc_63 <= th_myfunc_63_7;
        end
        th_myfunc_63_9: begin
          th_myfunc_63 <= th_myfunc_63_10;
        end
        th_myfunc_63_10: begin
          $display("Thread %d count = %d", _th_myfunc_63_tid_514, count);
          th_myfunc_63 <= th_myfunc_63_11;
        end
        th_myfunc_63_11: begin
          th_myfunc_63 <= th_myfunc_63_12;
        end
        th_myfunc_63_12: begin
          $display("Thread %d Unlock", _th_myfunc_63_tid_514);
          th_myfunc_63 <= th_myfunc_63_13;
        end
        th_myfunc_63_13: begin
          if((th_blink == 19) && (_th_blink_tid_260 == 63)) begin
            _th_myfunc_63_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_260 == 63)) begin
            th_myfunc_63 <= th_myfunc_63_init;
          end 
        end
      endcase
    end
  end


endmodule

