

module top
(
  input clk,
  input btnCpuReset,
  input btnC,
  input btnU,
  input btnL,
  input btnR,
  input btnD,
  input [16-1:0] sw,
  output [16-1:0] led
);

  wire new_CLK;
  assign new_CLK = clk;
  reg RST_X;
  reg RST;

  always @(posedge clk) begin
    RST_X <= btnCpuReset;
    RST <= !RST_X;
  end


  blinkled
  inst_blinkled
  (
    .CLK(new_CLK),
    .RST(RST),
    .btnC(btnC),
    .btnU(btnU),
    .btnL(btnL),
    .btnR(btnR),
    .btnD(btnD),
    .sw(sw),
    .led(led)
  );


endmodule



module blinkled
(
  input CLK,
  input RST,
  input btnC,
  input btnU,
  input btnL,
  input btnR,
  input btnD,
  input [16-1:0] sw,
  output [16-1:0] led
);

  reg [15-1:0] count;
  reg done;
  assign led = { done, count };
  reg _mymutex_lock_reg;
  reg [32-1:0] _mymutex_lock_id;
  reg [64-1:0] _th_myfunc_start;
  reg [32-1:0] th_blink;
  localparam th_blink_init = 0;
  reg signed [32-1:0] _th_blink_polarity_323;
  reg signed [32-1:0] _th_blink_tid_324;
  reg [32-1:0] th_myfunc_0;
  localparam th_myfunc_0_init = 0;
  reg [32-1:0] th_myfunc_1;
  localparam th_myfunc_1_init = 0;
  reg [32-1:0] th_myfunc_2;
  localparam th_myfunc_2_init = 0;
  reg [32-1:0] th_myfunc_3;
  localparam th_myfunc_3_init = 0;
  reg [32-1:0] th_myfunc_4;
  localparam th_myfunc_4_init = 0;
  reg [32-1:0] th_myfunc_5;
  localparam th_myfunc_5_init = 0;
  reg [32-1:0] th_myfunc_6;
  localparam th_myfunc_6_init = 0;
  reg [32-1:0] th_myfunc_7;
  localparam th_myfunc_7_init = 0;
  reg [32-1:0] th_myfunc_8;
  localparam th_myfunc_8_init = 0;
  reg [32-1:0] th_myfunc_9;
  localparam th_myfunc_9_init = 0;
  reg [32-1:0] th_myfunc_10;
  localparam th_myfunc_10_init = 0;
  reg [32-1:0] th_myfunc_11;
  localparam th_myfunc_11_init = 0;
  reg [32-1:0] th_myfunc_12;
  localparam th_myfunc_12_init = 0;
  reg [32-1:0] th_myfunc_13;
  localparam th_myfunc_13_init = 0;
  reg [32-1:0] th_myfunc_14;
  localparam th_myfunc_14_init = 0;
  reg [32-1:0] th_myfunc_15;
  localparam th_myfunc_15_init = 0;
  reg [32-1:0] th_myfunc_16;
  localparam th_myfunc_16_init = 0;
  reg [32-1:0] th_myfunc_17;
  localparam th_myfunc_17_init = 0;
  reg [32-1:0] th_myfunc_18;
  localparam th_myfunc_18_init = 0;
  reg [32-1:0] th_myfunc_19;
  localparam th_myfunc_19_init = 0;
  reg [32-1:0] th_myfunc_20;
  localparam th_myfunc_20_init = 0;
  reg [32-1:0] th_myfunc_21;
  localparam th_myfunc_21_init = 0;
  reg [32-1:0] th_myfunc_22;
  localparam th_myfunc_22_init = 0;
  reg [32-1:0] th_myfunc_23;
  localparam th_myfunc_23_init = 0;
  reg [32-1:0] th_myfunc_24;
  localparam th_myfunc_24_init = 0;
  reg [32-1:0] th_myfunc_25;
  localparam th_myfunc_25_init = 0;
  reg [32-1:0] th_myfunc_26;
  localparam th_myfunc_26_init = 0;
  reg [32-1:0] th_myfunc_27;
  localparam th_myfunc_27_init = 0;
  reg [32-1:0] th_myfunc_28;
  localparam th_myfunc_28_init = 0;
  reg [32-1:0] th_myfunc_29;
  localparam th_myfunc_29_init = 0;
  reg [32-1:0] th_myfunc_30;
  localparam th_myfunc_30_init = 0;
  reg [32-1:0] th_myfunc_31;
  localparam th_myfunc_31_init = 0;
  reg [32-1:0] th_myfunc_32;
  localparam th_myfunc_32_init = 0;
  reg [32-1:0] th_myfunc_33;
  localparam th_myfunc_33_init = 0;
  reg [32-1:0] th_myfunc_34;
  localparam th_myfunc_34_init = 0;
  reg [32-1:0] th_myfunc_35;
  localparam th_myfunc_35_init = 0;
  reg [32-1:0] th_myfunc_36;
  localparam th_myfunc_36_init = 0;
  reg [32-1:0] th_myfunc_37;
  localparam th_myfunc_37_init = 0;
  reg [32-1:0] th_myfunc_38;
  localparam th_myfunc_38_init = 0;
  reg [32-1:0] th_myfunc_39;
  localparam th_myfunc_39_init = 0;
  reg [32-1:0] th_myfunc_40;
  localparam th_myfunc_40_init = 0;
  reg [32-1:0] th_myfunc_41;
  localparam th_myfunc_41_init = 0;
  reg [32-1:0] th_myfunc_42;
  localparam th_myfunc_42_init = 0;
  reg [32-1:0] th_myfunc_43;
  localparam th_myfunc_43_init = 0;
  reg [32-1:0] th_myfunc_44;
  localparam th_myfunc_44_init = 0;
  reg [32-1:0] th_myfunc_45;
  localparam th_myfunc_45_init = 0;
  reg [32-1:0] th_myfunc_46;
  localparam th_myfunc_46_init = 0;
  reg [32-1:0] th_myfunc_47;
  localparam th_myfunc_47_init = 0;
  reg [32-1:0] th_myfunc_48;
  localparam th_myfunc_48_init = 0;
  reg [32-1:0] th_myfunc_49;
  localparam th_myfunc_49_init = 0;
  reg [32-1:0] th_myfunc_50;
  localparam th_myfunc_50_init = 0;
  reg [32-1:0] th_myfunc_51;
  localparam th_myfunc_51_init = 0;
  reg [32-1:0] th_myfunc_52;
  localparam th_myfunc_52_init = 0;
  reg [32-1:0] th_myfunc_53;
  localparam th_myfunc_53_init = 0;
  reg [32-1:0] th_myfunc_54;
  localparam th_myfunc_54_init = 0;
  reg [32-1:0] th_myfunc_55;
  localparam th_myfunc_55_init = 0;
  reg [32-1:0] th_myfunc_56;
  localparam th_myfunc_56_init = 0;
  reg [32-1:0] th_myfunc_57;
  localparam th_myfunc_57_init = 0;
  reg [32-1:0] th_myfunc_58;
  localparam th_myfunc_58_init = 0;
  reg [32-1:0] th_myfunc_59;
  localparam th_myfunc_59_init = 0;
  reg [32-1:0] th_myfunc_60;
  localparam th_myfunc_60_init = 0;
  reg [32-1:0] th_myfunc_61;
  localparam th_myfunc_61_init = 0;
  reg [32-1:0] th_myfunc_62;
  localparam th_myfunc_62_init = 0;
  reg [32-1:0] th_myfunc_63;
  localparam th_myfunc_63_init = 0;
  reg _th_myfunc_0_called;
  reg signed [32-1:0] _th_myfunc_0_tid_325;
  reg signed [32-1:0] _th_myfunc_0_tid_326;
  reg signed [32-1:0] _th_myfunc_0_time_327;
  reg signed [32-1:0] _th_myfunc_0_i_328;
  reg signed [32-1:0] _th_myfunc_0___329;
  reg _th_myfunc_1_called;
  reg signed [32-1:0] _th_myfunc_1_tid_330;
  reg signed [32-1:0] _th_myfunc_1_tid_331;
  reg signed [32-1:0] _th_myfunc_1_time_332;
  reg signed [32-1:0] _th_myfunc_1_i_333;
  reg signed [32-1:0] _th_myfunc_1___334;
  reg _th_myfunc_2_called;
  reg signed [32-1:0] _th_myfunc_2_tid_335;
  reg signed [32-1:0] _th_myfunc_2_tid_336;
  reg signed [32-1:0] _th_myfunc_2_time_337;
  reg signed [32-1:0] _th_myfunc_2_i_338;
  reg signed [32-1:0] _th_myfunc_2___339;
  reg _th_myfunc_3_called;
  reg signed [32-1:0] _th_myfunc_3_tid_340;
  reg signed [32-1:0] _th_myfunc_3_tid_341;
  reg signed [32-1:0] _th_myfunc_3_time_342;
  reg signed [32-1:0] _th_myfunc_3_i_343;
  reg signed [32-1:0] _th_myfunc_3___344;
  reg _th_myfunc_4_called;
  reg signed [32-1:0] _th_myfunc_4_tid_345;
  reg signed [32-1:0] _th_myfunc_4_tid_346;
  reg signed [32-1:0] _th_myfunc_4_time_347;
  reg signed [32-1:0] _th_myfunc_4_i_348;
  reg signed [32-1:0] _th_myfunc_4___349;
  reg _th_myfunc_5_called;
  reg signed [32-1:0] _th_myfunc_5_tid_350;
  reg signed [32-1:0] _th_myfunc_5_tid_351;
  reg signed [32-1:0] _th_myfunc_5_time_352;
  reg signed [32-1:0] _th_myfunc_5_i_353;
  reg signed [32-1:0] _th_myfunc_5___354;
  reg _th_myfunc_6_called;
  reg signed [32-1:0] _th_myfunc_6_tid_355;
  reg signed [32-1:0] _th_myfunc_6_tid_356;
  reg signed [32-1:0] _th_myfunc_6_time_357;
  reg signed [32-1:0] _th_myfunc_6_i_358;
  reg signed [32-1:0] _th_myfunc_6___359;
  reg _th_myfunc_7_called;
  reg signed [32-1:0] _th_myfunc_7_tid_360;
  reg signed [32-1:0] _th_myfunc_7_tid_361;
  reg signed [32-1:0] _th_myfunc_7_time_362;
  reg signed [32-1:0] _th_myfunc_7_i_363;
  reg signed [32-1:0] _th_myfunc_7___364;
  reg _th_myfunc_8_called;
  reg signed [32-1:0] _th_myfunc_8_tid_365;
  reg signed [32-1:0] _th_myfunc_8_tid_366;
  reg signed [32-1:0] _th_myfunc_8_time_367;
  reg signed [32-1:0] _th_myfunc_8_i_368;
  reg signed [32-1:0] _th_myfunc_8___369;
  reg _th_myfunc_9_called;
  reg signed [32-1:0] _th_myfunc_9_tid_370;
  reg signed [32-1:0] _th_myfunc_9_tid_371;
  reg signed [32-1:0] _th_myfunc_9_time_372;
  reg signed [32-1:0] _th_myfunc_9_i_373;
  reg signed [32-1:0] _th_myfunc_9___374;
  reg _th_myfunc_10_called;
  reg signed [32-1:0] _th_myfunc_10_tid_375;
  reg signed [32-1:0] _th_myfunc_10_tid_376;
  reg signed [32-1:0] _th_myfunc_10_time_377;
  reg signed [32-1:0] _th_myfunc_10_i_378;
  reg signed [32-1:0] _th_myfunc_10___379;
  reg _th_myfunc_11_called;
  reg signed [32-1:0] _th_myfunc_11_tid_380;
  reg signed [32-1:0] _th_myfunc_11_tid_381;
  reg signed [32-1:0] _th_myfunc_11_time_382;
  reg signed [32-1:0] _th_myfunc_11_i_383;
  reg signed [32-1:0] _th_myfunc_11___384;
  reg _th_myfunc_12_called;
  reg signed [32-1:0] _th_myfunc_12_tid_385;
  reg signed [32-1:0] _th_myfunc_12_tid_386;
  reg signed [32-1:0] _th_myfunc_12_time_387;
  reg signed [32-1:0] _th_myfunc_12_i_388;
  reg signed [32-1:0] _th_myfunc_12___389;
  reg _th_myfunc_13_called;
  reg signed [32-1:0] _th_myfunc_13_tid_390;
  reg signed [32-1:0] _th_myfunc_13_tid_391;
  reg signed [32-1:0] _th_myfunc_13_time_392;
  reg signed [32-1:0] _th_myfunc_13_i_393;
  reg signed [32-1:0] _th_myfunc_13___394;
  reg _th_myfunc_14_called;
  reg signed [32-1:0] _th_myfunc_14_tid_395;
  reg signed [32-1:0] _th_myfunc_14_tid_396;
  reg signed [32-1:0] _th_myfunc_14_time_397;
  reg signed [32-1:0] _th_myfunc_14_i_398;
  reg signed [32-1:0] _th_myfunc_14___399;
  reg _th_myfunc_15_called;
  reg signed [32-1:0] _th_myfunc_15_tid_400;
  reg signed [32-1:0] _th_myfunc_15_tid_401;
  reg signed [32-1:0] _th_myfunc_15_time_402;
  reg signed [32-1:0] _th_myfunc_15_i_403;
  reg signed [32-1:0] _th_myfunc_15___404;
  reg _th_myfunc_16_called;
  reg signed [32-1:0] _th_myfunc_16_tid_405;
  reg signed [32-1:0] _th_myfunc_16_tid_406;
  reg signed [32-1:0] _th_myfunc_16_time_407;
  reg signed [32-1:0] _th_myfunc_16_i_408;
  reg signed [32-1:0] _th_myfunc_16___409;
  reg _th_myfunc_17_called;
  reg signed [32-1:0] _th_myfunc_17_tid_410;
  reg signed [32-1:0] _th_myfunc_17_tid_411;
  reg signed [32-1:0] _th_myfunc_17_time_412;
  reg signed [32-1:0] _th_myfunc_17_i_413;
  reg signed [32-1:0] _th_myfunc_17___414;
  reg _th_myfunc_18_called;
  reg signed [32-1:0] _th_myfunc_18_tid_415;
  reg signed [32-1:0] _th_myfunc_18_tid_416;
  reg signed [32-1:0] _th_myfunc_18_time_417;
  reg signed [32-1:0] _th_myfunc_18_i_418;
  reg signed [32-1:0] _th_myfunc_18___419;
  reg _th_myfunc_19_called;
  reg signed [32-1:0] _th_myfunc_19_tid_420;
  reg signed [32-1:0] _th_myfunc_19_tid_421;
  reg signed [32-1:0] _th_myfunc_19_time_422;
  reg signed [32-1:0] _th_myfunc_19_i_423;
  reg signed [32-1:0] _th_myfunc_19___424;
  reg _th_myfunc_20_called;
  reg signed [32-1:0] _th_myfunc_20_tid_425;
  reg signed [32-1:0] _th_myfunc_20_tid_426;
  reg signed [32-1:0] _th_myfunc_20_time_427;
  reg signed [32-1:0] _th_myfunc_20_i_428;
  reg signed [32-1:0] _th_myfunc_20___429;
  reg _th_myfunc_21_called;
  reg signed [32-1:0] _th_myfunc_21_tid_430;
  reg signed [32-1:0] _th_myfunc_21_tid_431;
  reg signed [32-1:0] _th_myfunc_21_time_432;
  reg signed [32-1:0] _th_myfunc_21_i_433;
  reg signed [32-1:0] _th_myfunc_21___434;
  reg _th_myfunc_22_called;
  reg signed [32-1:0] _th_myfunc_22_tid_435;
  reg signed [32-1:0] _th_myfunc_22_tid_436;
  reg signed [32-1:0] _th_myfunc_22_time_437;
  reg signed [32-1:0] _th_myfunc_22_i_438;
  reg signed [32-1:0] _th_myfunc_22___439;
  reg _th_myfunc_23_called;
  reg signed [32-1:0] _th_myfunc_23_tid_440;
  reg signed [32-1:0] _th_myfunc_23_tid_441;
  reg signed [32-1:0] _th_myfunc_23_time_442;
  reg signed [32-1:0] _th_myfunc_23_i_443;
  reg signed [32-1:0] _th_myfunc_23___444;
  reg _th_myfunc_24_called;
  reg signed [32-1:0] _th_myfunc_24_tid_445;
  reg signed [32-1:0] _th_myfunc_24_tid_446;
  reg signed [32-1:0] _th_myfunc_24_time_447;
  reg signed [32-1:0] _th_myfunc_24_i_448;
  reg signed [32-1:0] _th_myfunc_24___449;
  reg _th_myfunc_25_called;
  reg signed [32-1:0] _th_myfunc_25_tid_450;
  reg signed [32-1:0] _th_myfunc_25_tid_451;
  reg signed [32-1:0] _th_myfunc_25_time_452;
  reg signed [32-1:0] _th_myfunc_25_i_453;
  reg signed [32-1:0] _th_myfunc_25___454;
  reg _th_myfunc_26_called;
  reg signed [32-1:0] _th_myfunc_26_tid_455;
  reg signed [32-1:0] _th_myfunc_26_tid_456;
  reg signed [32-1:0] _th_myfunc_26_time_457;
  reg signed [32-1:0] _th_myfunc_26_i_458;
  reg signed [32-1:0] _th_myfunc_26___459;
  reg _th_myfunc_27_called;
  reg signed [32-1:0] _th_myfunc_27_tid_460;
  reg signed [32-1:0] _th_myfunc_27_tid_461;
  reg signed [32-1:0] _th_myfunc_27_time_462;
  reg signed [32-1:0] _th_myfunc_27_i_463;
  reg signed [32-1:0] _th_myfunc_27___464;
  reg _th_myfunc_28_called;
  reg signed [32-1:0] _th_myfunc_28_tid_465;
  reg signed [32-1:0] _th_myfunc_28_tid_466;
  reg signed [32-1:0] _th_myfunc_28_time_467;
  reg signed [32-1:0] _th_myfunc_28_i_468;
  reg signed [32-1:0] _th_myfunc_28___469;
  reg _th_myfunc_29_called;
  reg signed [32-1:0] _th_myfunc_29_tid_470;
  reg signed [32-1:0] _th_myfunc_29_tid_471;
  reg signed [32-1:0] _th_myfunc_29_time_472;
  reg signed [32-1:0] _th_myfunc_29_i_473;
  reg signed [32-1:0] _th_myfunc_29___474;
  reg _th_myfunc_30_called;
  reg signed [32-1:0] _th_myfunc_30_tid_475;
  reg signed [32-1:0] _th_myfunc_30_tid_476;
  reg signed [32-1:0] _th_myfunc_30_time_477;
  reg signed [32-1:0] _th_myfunc_30_i_478;
  reg signed [32-1:0] _th_myfunc_30___479;
  reg _th_myfunc_31_called;
  reg signed [32-1:0] _th_myfunc_31_tid_480;
  reg signed [32-1:0] _th_myfunc_31_tid_481;
  reg signed [32-1:0] _th_myfunc_31_time_482;
  reg signed [32-1:0] _th_myfunc_31_i_483;
  reg signed [32-1:0] _th_myfunc_31___484;
  reg _th_myfunc_32_called;
  reg signed [32-1:0] _th_myfunc_32_tid_485;
  reg signed [32-1:0] _th_myfunc_32_tid_486;
  reg signed [32-1:0] _th_myfunc_32_time_487;
  reg signed [32-1:0] _th_myfunc_32_i_488;
  reg signed [32-1:0] _th_myfunc_32___489;
  reg _th_myfunc_33_called;
  reg signed [32-1:0] _th_myfunc_33_tid_490;
  reg signed [32-1:0] _th_myfunc_33_tid_491;
  reg signed [32-1:0] _th_myfunc_33_time_492;
  reg signed [32-1:0] _th_myfunc_33_i_493;
  reg signed [32-1:0] _th_myfunc_33___494;
  reg _th_myfunc_34_called;
  reg signed [32-1:0] _th_myfunc_34_tid_495;
  reg signed [32-1:0] _th_myfunc_34_tid_496;
  reg signed [32-1:0] _th_myfunc_34_time_497;
  reg signed [32-1:0] _th_myfunc_34_i_498;
  reg signed [32-1:0] _th_myfunc_34___499;
  reg _th_myfunc_35_called;
  reg signed [32-1:0] _th_myfunc_35_tid_500;
  reg signed [32-1:0] _th_myfunc_35_tid_501;
  reg signed [32-1:0] _th_myfunc_35_time_502;
  reg signed [32-1:0] _th_myfunc_35_i_503;
  reg signed [32-1:0] _th_myfunc_35___504;
  reg _th_myfunc_36_called;
  reg signed [32-1:0] _th_myfunc_36_tid_505;
  reg signed [32-1:0] _th_myfunc_36_tid_506;
  reg signed [32-1:0] _th_myfunc_36_time_507;
  reg signed [32-1:0] _th_myfunc_36_i_508;
  reg signed [32-1:0] _th_myfunc_36___509;
  reg _th_myfunc_37_called;
  reg signed [32-1:0] _th_myfunc_37_tid_510;
  reg signed [32-1:0] _th_myfunc_37_tid_511;
  reg signed [32-1:0] _th_myfunc_37_time_512;
  reg signed [32-1:0] _th_myfunc_37_i_513;
  reg signed [32-1:0] _th_myfunc_37___514;
  reg _th_myfunc_38_called;
  reg signed [32-1:0] _th_myfunc_38_tid_515;
  reg signed [32-1:0] _th_myfunc_38_tid_516;
  reg signed [32-1:0] _th_myfunc_38_time_517;
  reg signed [32-1:0] _th_myfunc_38_i_518;
  reg signed [32-1:0] _th_myfunc_38___519;
  reg _th_myfunc_39_called;
  reg signed [32-1:0] _th_myfunc_39_tid_520;
  reg signed [32-1:0] _th_myfunc_39_tid_521;
  reg signed [32-1:0] _th_myfunc_39_time_522;
  reg signed [32-1:0] _th_myfunc_39_i_523;
  reg signed [32-1:0] _th_myfunc_39___524;
  reg _th_myfunc_40_called;
  reg signed [32-1:0] _th_myfunc_40_tid_525;
  reg signed [32-1:0] _th_myfunc_40_tid_526;
  reg signed [32-1:0] _th_myfunc_40_time_527;
  reg signed [32-1:0] _th_myfunc_40_i_528;
  reg signed [32-1:0] _th_myfunc_40___529;
  reg _th_myfunc_41_called;
  reg signed [32-1:0] _th_myfunc_41_tid_530;
  reg signed [32-1:0] _th_myfunc_41_tid_531;
  reg signed [32-1:0] _th_myfunc_41_time_532;
  reg signed [32-1:0] _th_myfunc_41_i_533;
  reg signed [32-1:0] _th_myfunc_41___534;
  reg _th_myfunc_42_called;
  reg signed [32-1:0] _th_myfunc_42_tid_535;
  reg signed [32-1:0] _th_myfunc_42_tid_536;
  reg signed [32-1:0] _th_myfunc_42_time_537;
  reg signed [32-1:0] _th_myfunc_42_i_538;
  reg signed [32-1:0] _th_myfunc_42___539;
  reg _th_myfunc_43_called;
  reg signed [32-1:0] _th_myfunc_43_tid_540;
  reg signed [32-1:0] _th_myfunc_43_tid_541;
  reg signed [32-1:0] _th_myfunc_43_time_542;
  reg signed [32-1:0] _th_myfunc_43_i_543;
  reg signed [32-1:0] _th_myfunc_43___544;
  reg _th_myfunc_44_called;
  reg signed [32-1:0] _th_myfunc_44_tid_545;
  reg signed [32-1:0] _th_myfunc_44_tid_546;
  reg signed [32-1:0] _th_myfunc_44_time_547;
  reg signed [32-1:0] _th_myfunc_44_i_548;
  reg signed [32-1:0] _th_myfunc_44___549;
  reg _th_myfunc_45_called;
  reg signed [32-1:0] _th_myfunc_45_tid_550;
  reg signed [32-1:0] _th_myfunc_45_tid_551;
  reg signed [32-1:0] _th_myfunc_45_time_552;
  reg signed [32-1:0] _th_myfunc_45_i_553;
  reg signed [32-1:0] _th_myfunc_45___554;
  reg _th_myfunc_46_called;
  reg signed [32-1:0] _th_myfunc_46_tid_555;
  reg signed [32-1:0] _th_myfunc_46_tid_556;
  reg signed [32-1:0] _th_myfunc_46_time_557;
  reg signed [32-1:0] _th_myfunc_46_i_558;
  reg signed [32-1:0] _th_myfunc_46___559;
  reg _th_myfunc_47_called;
  reg signed [32-1:0] _th_myfunc_47_tid_560;
  reg signed [32-1:0] _th_myfunc_47_tid_561;
  reg signed [32-1:0] _th_myfunc_47_time_562;
  reg signed [32-1:0] _th_myfunc_47_i_563;
  reg signed [32-1:0] _th_myfunc_47___564;
  reg _th_myfunc_48_called;
  reg signed [32-1:0] _th_myfunc_48_tid_565;
  reg signed [32-1:0] _th_myfunc_48_tid_566;
  reg signed [32-1:0] _th_myfunc_48_time_567;
  reg signed [32-1:0] _th_myfunc_48_i_568;
  reg signed [32-1:0] _th_myfunc_48___569;
  reg _th_myfunc_49_called;
  reg signed [32-1:0] _th_myfunc_49_tid_570;
  reg signed [32-1:0] _th_myfunc_49_tid_571;
  reg signed [32-1:0] _th_myfunc_49_time_572;
  reg signed [32-1:0] _th_myfunc_49_i_573;
  reg signed [32-1:0] _th_myfunc_49___574;
  reg _th_myfunc_50_called;
  reg signed [32-1:0] _th_myfunc_50_tid_575;
  reg signed [32-1:0] _th_myfunc_50_tid_576;
  reg signed [32-1:0] _th_myfunc_50_time_577;
  reg signed [32-1:0] _th_myfunc_50_i_578;
  reg signed [32-1:0] _th_myfunc_50___579;
  reg _th_myfunc_51_called;
  reg signed [32-1:0] _th_myfunc_51_tid_580;
  reg signed [32-1:0] _th_myfunc_51_tid_581;
  reg signed [32-1:0] _th_myfunc_51_time_582;
  reg signed [32-1:0] _th_myfunc_51_i_583;
  reg signed [32-1:0] _th_myfunc_51___584;
  reg _th_myfunc_52_called;
  reg signed [32-1:0] _th_myfunc_52_tid_585;
  reg signed [32-1:0] _th_myfunc_52_tid_586;
  reg signed [32-1:0] _th_myfunc_52_time_587;
  reg signed [32-1:0] _th_myfunc_52_i_588;
  reg signed [32-1:0] _th_myfunc_52___589;
  reg _th_myfunc_53_called;
  reg signed [32-1:0] _th_myfunc_53_tid_590;
  reg signed [32-1:0] _th_myfunc_53_tid_591;
  reg signed [32-1:0] _th_myfunc_53_time_592;
  reg signed [32-1:0] _th_myfunc_53_i_593;
  reg signed [32-1:0] _th_myfunc_53___594;
  reg _th_myfunc_54_called;
  reg signed [32-1:0] _th_myfunc_54_tid_595;
  reg signed [32-1:0] _th_myfunc_54_tid_596;
  reg signed [32-1:0] _th_myfunc_54_time_597;
  reg signed [32-1:0] _th_myfunc_54_i_598;
  reg signed [32-1:0] _th_myfunc_54___599;
  reg _th_myfunc_55_called;
  reg signed [32-1:0] _th_myfunc_55_tid_600;
  reg signed [32-1:0] _th_myfunc_55_tid_601;
  reg signed [32-1:0] _th_myfunc_55_time_602;
  reg signed [32-1:0] _th_myfunc_55_i_603;
  reg signed [32-1:0] _th_myfunc_55___604;
  reg _th_myfunc_56_called;
  reg signed [32-1:0] _th_myfunc_56_tid_605;
  reg signed [32-1:0] _th_myfunc_56_tid_606;
  reg signed [32-1:0] _th_myfunc_56_time_607;
  reg signed [32-1:0] _th_myfunc_56_i_608;
  reg signed [32-1:0] _th_myfunc_56___609;
  reg _th_myfunc_57_called;
  reg signed [32-1:0] _th_myfunc_57_tid_610;
  reg signed [32-1:0] _th_myfunc_57_tid_611;
  reg signed [32-1:0] _th_myfunc_57_time_612;
  reg signed [32-1:0] _th_myfunc_57_i_613;
  reg signed [32-1:0] _th_myfunc_57___614;
  reg _th_myfunc_58_called;
  reg signed [32-1:0] _th_myfunc_58_tid_615;
  reg signed [32-1:0] _th_myfunc_58_tid_616;
  reg signed [32-1:0] _th_myfunc_58_time_617;
  reg signed [32-1:0] _th_myfunc_58_i_618;
  reg signed [32-1:0] _th_myfunc_58___619;
  reg _th_myfunc_59_called;
  reg signed [32-1:0] _th_myfunc_59_tid_620;
  reg signed [32-1:0] _th_myfunc_59_tid_621;
  reg signed [32-1:0] _th_myfunc_59_time_622;
  reg signed [32-1:0] _th_myfunc_59_i_623;
  reg signed [32-1:0] _th_myfunc_59___624;
  reg _th_myfunc_60_called;
  reg signed [32-1:0] _th_myfunc_60_tid_625;
  reg signed [32-1:0] _th_myfunc_60_tid_626;
  reg signed [32-1:0] _th_myfunc_60_time_627;
  reg signed [32-1:0] _th_myfunc_60_i_628;
  reg signed [32-1:0] _th_myfunc_60___629;
  reg _th_myfunc_61_called;
  reg signed [32-1:0] _th_myfunc_61_tid_630;
  reg signed [32-1:0] _th_myfunc_61_tid_631;
  reg signed [32-1:0] _th_myfunc_61_time_632;
  reg signed [32-1:0] _th_myfunc_61_i_633;
  reg signed [32-1:0] _th_myfunc_61___634;
  reg _th_myfunc_62_called;
  reg signed [32-1:0] _th_myfunc_62_tid_635;
  reg signed [32-1:0] _th_myfunc_62_tid_636;
  reg signed [32-1:0] _th_myfunc_62_time_637;
  reg signed [32-1:0] _th_myfunc_62_i_638;
  reg signed [32-1:0] _th_myfunc_62___639;
  reg _th_myfunc_63_called;
  reg signed [32-1:0] _th_myfunc_63_tid_640;
  reg signed [32-1:0] _th_myfunc_63_tid_641;
  reg signed [32-1:0] _th_myfunc_63_time_642;
  reg signed [32-1:0] _th_myfunc_63_i_643;
  reg signed [32-1:0] _th_myfunc_63___644;

  always @(posedge CLK) begin
    if(RST) begin
      _mymutex_lock_reg <= 0;
      _mymutex_lock_id <= 0;
    end else begin
      if((th_myfunc_0 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 0;
      end 
      if((th_myfunc_0 == 14) && (_mymutex_lock_id == 0)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_1 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 1;
      end 
      if((th_myfunc_1 == 14) && (_mymutex_lock_id == 1)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_2 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 2;
      end 
      if((th_myfunc_2 == 14) && (_mymutex_lock_id == 2)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_3 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 3;
      end 
      if((th_myfunc_3 == 14) && (_mymutex_lock_id == 3)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_4 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 4;
      end 
      if((th_myfunc_4 == 14) && (_mymutex_lock_id == 4)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_5 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 5;
      end 
      if((th_myfunc_5 == 14) && (_mymutex_lock_id == 5)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_6 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 6;
      end 
      if((th_myfunc_6 == 14) && (_mymutex_lock_id == 6)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_7 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 7;
      end 
      if((th_myfunc_7 == 14) && (_mymutex_lock_id == 7)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_8 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 8;
      end 
      if((th_myfunc_8 == 14) && (_mymutex_lock_id == 8)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_9 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 9;
      end 
      if((th_myfunc_9 == 14) && (_mymutex_lock_id == 9)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_10 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 10;
      end 
      if((th_myfunc_10 == 14) && (_mymutex_lock_id == 10)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_11 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 11;
      end 
      if((th_myfunc_11 == 14) && (_mymutex_lock_id == 11)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_12 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 12;
      end 
      if((th_myfunc_12 == 14) && (_mymutex_lock_id == 12)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_13 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 13;
      end 
      if((th_myfunc_13 == 14) && (_mymutex_lock_id == 13)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_14 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 14;
      end 
      if((th_myfunc_14 == 14) && (_mymutex_lock_id == 14)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_15 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 15;
      end 
      if((th_myfunc_15 == 14) && (_mymutex_lock_id == 15)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_16 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 16;
      end 
      if((th_myfunc_16 == 14) && (_mymutex_lock_id == 16)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_17 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 17;
      end 
      if((th_myfunc_17 == 14) && (_mymutex_lock_id == 17)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_18 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 18;
      end 
      if((th_myfunc_18 == 14) && (_mymutex_lock_id == 18)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_19 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 19;
      end 
      if((th_myfunc_19 == 14) && (_mymutex_lock_id == 19)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_20 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 20;
      end 
      if((th_myfunc_20 == 14) && (_mymutex_lock_id == 20)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_21 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 21;
      end 
      if((th_myfunc_21 == 14) && (_mymutex_lock_id == 21)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_22 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 22;
      end 
      if((th_myfunc_22 == 14) && (_mymutex_lock_id == 22)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_23 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 23;
      end 
      if((th_myfunc_23 == 14) && (_mymutex_lock_id == 23)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_24 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 24;
      end 
      if((th_myfunc_24 == 14) && (_mymutex_lock_id == 24)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_25 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 25;
      end 
      if((th_myfunc_25 == 14) && (_mymutex_lock_id == 25)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_26 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 26;
      end 
      if((th_myfunc_26 == 14) && (_mymutex_lock_id == 26)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_27 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 27;
      end 
      if((th_myfunc_27 == 14) && (_mymutex_lock_id == 27)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_28 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 28;
      end 
      if((th_myfunc_28 == 14) && (_mymutex_lock_id == 28)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_29 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 29;
      end 
      if((th_myfunc_29 == 14) && (_mymutex_lock_id == 29)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_30 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 30;
      end 
      if((th_myfunc_30 == 14) && (_mymutex_lock_id == 30)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_31 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 31;
      end 
      if((th_myfunc_31 == 14) && (_mymutex_lock_id == 31)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_32 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 32;
      end 
      if((th_myfunc_32 == 14) && (_mymutex_lock_id == 32)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_33 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 33;
      end 
      if((th_myfunc_33 == 14) && (_mymutex_lock_id == 33)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_34 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 34;
      end 
      if((th_myfunc_34 == 14) && (_mymutex_lock_id == 34)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_35 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 35;
      end 
      if((th_myfunc_35 == 14) && (_mymutex_lock_id == 35)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_36 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 36;
      end 
      if((th_myfunc_36 == 14) && (_mymutex_lock_id == 36)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_37 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 37;
      end 
      if((th_myfunc_37 == 14) && (_mymutex_lock_id == 37)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_38 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 38;
      end 
      if((th_myfunc_38 == 14) && (_mymutex_lock_id == 38)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_39 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 39;
      end 
      if((th_myfunc_39 == 14) && (_mymutex_lock_id == 39)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_40 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 40;
      end 
      if((th_myfunc_40 == 14) && (_mymutex_lock_id == 40)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_41 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 41;
      end 
      if((th_myfunc_41 == 14) && (_mymutex_lock_id == 41)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_42 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 42;
      end 
      if((th_myfunc_42 == 14) && (_mymutex_lock_id == 42)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_43 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 43;
      end 
      if((th_myfunc_43 == 14) && (_mymutex_lock_id == 43)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_44 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 44;
      end 
      if((th_myfunc_44 == 14) && (_mymutex_lock_id == 44)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_45 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 45;
      end 
      if((th_myfunc_45 == 14) && (_mymutex_lock_id == 45)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_46 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 46;
      end 
      if((th_myfunc_46 == 14) && (_mymutex_lock_id == 46)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_47 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 47;
      end 
      if((th_myfunc_47 == 14) && (_mymutex_lock_id == 47)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_48 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 48;
      end 
      if((th_myfunc_48 == 14) && (_mymutex_lock_id == 48)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_49 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 49;
      end 
      if((th_myfunc_49 == 14) && (_mymutex_lock_id == 49)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_50 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 50;
      end 
      if((th_myfunc_50 == 14) && (_mymutex_lock_id == 50)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_51 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 51;
      end 
      if((th_myfunc_51 == 14) && (_mymutex_lock_id == 51)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_52 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 52;
      end 
      if((th_myfunc_52 == 14) && (_mymutex_lock_id == 52)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_53 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 53;
      end 
      if((th_myfunc_53 == 14) && (_mymutex_lock_id == 53)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_54 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 54;
      end 
      if((th_myfunc_54 == 14) && (_mymutex_lock_id == 54)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_55 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 55;
      end 
      if((th_myfunc_55 == 14) && (_mymutex_lock_id == 55)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_56 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 56;
      end 
      if((th_myfunc_56 == 14) && (_mymutex_lock_id == 56)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_57 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 57;
      end 
      if((th_myfunc_57 == 14) && (_mymutex_lock_id == 57)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_58 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 58;
      end 
      if((th_myfunc_58 == 14) && (_mymutex_lock_id == 58)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_59 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 59;
      end 
      if((th_myfunc_59 == 14) && (_mymutex_lock_id == 59)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_60 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 60;
      end 
      if((th_myfunc_60 == 14) && (_mymutex_lock_id == 60)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_61 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 61;
      end 
      if((th_myfunc_61 == 14) && (_mymutex_lock_id == 61)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_62 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 62;
      end 
      if((th_myfunc_62 == 14) && (_mymutex_lock_id == 62)) begin
        _mymutex_lock_reg <= 0;
      end 
      if((th_myfunc_63 == 2) && !_mymutex_lock_reg) begin
        _mymutex_lock_reg <= 1;
        _mymutex_lock_id <= 63;
      end 
      if((th_myfunc_63 == 14) && (_mymutex_lock_id == 63)) begin
        _mymutex_lock_reg <= 0;
      end 
    end
  end

  localparam th_blink_1 = 1;
  localparam th_blink_2 = 2;
  localparam th_blink_3 = 3;
  localparam th_blink_4 = 4;
  localparam th_blink_5 = 5;
  localparam th_blink_6 = 6;
  localparam th_blink_7 = 7;
  localparam th_blink_8 = 8;
  localparam th_blink_9 = 9;
  localparam th_blink_10 = 10;
  localparam th_blink_11 = 11;
  localparam th_blink_12 = 12;
  localparam th_blink_13 = 13;
  localparam th_blink_14 = 14;
  localparam th_blink_15 = 15;
  localparam th_blink_16 = 16;
  localparam th_blink_17 = 17;
  localparam th_blink_18 = 18;
  localparam th_blink_19 = 19;
  localparam th_blink_20 = 20;
  localparam th_blink_21 = 21;
  localparam th_blink_22 = 22;

  always @(posedge CLK) begin
    if(RST) begin
      th_blink <= th_blink_init;
      done <= 0;
      _th_blink_polarity_323 <= 0;
      _th_blink_tid_324 <= 0;
      _th_myfunc_start[_th_blink_tid_324] <= (0 >> _th_blink_tid_324) & 1'd1;
    end else begin
      case(th_blink)
        th_blink_init: begin
          th_blink <= th_blink_1;
        end
        th_blink_1: begin
          th_blink <= th_blink_2;
        end
        th_blink_2: begin
          if(1) begin
            th_blink <= th_blink_3;
          end else begin
            th_blink <= th_blink_22;
          end
        end
        th_blink_3: begin
          done <= 0;
          th_blink <= th_blink_4;
        end
        th_blink_4: begin
          _th_blink_polarity_323 <= 1;
          th_blink <= th_blink_5;
        end
        th_blink_5: begin
          if(btnC != _th_blink_polarity_323) begin
            th_blink <= th_blink_6;
          end else begin
            th_blink <= th_blink_7;
          end
        end
        th_blink_6: begin
          th_blink <= th_blink_5;
        end
        th_blink_7: begin
          _th_blink_tid_324 <= 0;
          th_blink <= th_blink_8;
        end
        th_blink_8: begin
          if(_th_blink_tid_324 < 64) begin
            th_blink <= th_blink_9;
          end else begin
            th_blink <= th_blink_13;
          end
        end
        th_blink_9: begin
          _th_myfunc_start[_th_blink_tid_324] <= 1;
          th_blink <= th_blink_10;
        end
        th_blink_10: begin
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
          th_blink <= th_blink_11;
        end
        th_blink_11: begin
          _th_myfunc_start[_th_blink_tid_324] <= 0;
          th_blink <= th_blink_12;
        end
        th_blink_12: begin
          _th_blink_tid_324 <= _th_blink_tid_324 + 1;
          th_blink <= th_blink_8;
        end
        th_blink_13: begin
          _th_blink_tid_324 <= 0;
          th_blink <= th_blink_14;
        end
        th_blink_14: begin
          if(_th_blink_tid_324 < 64) begin
            th_blink <= th_blink_15;
          end else begin
            th_blink <= th_blink_17;
          end
        end
        th_blink_15: begin
          if((_th_blink_tid_324 == 0)? th_myfunc_0 == 16 : 
          (_th_blink_tid_324 == 1)? th_myfunc_1 == 16 : 
          (_th_blink_tid_324 == 2)? th_myfunc_2 == 16 : 
          (_th_blink_tid_324 == 3)? th_myfunc_3 == 16 : 
          (_th_blink_tid_324 == 4)? th_myfunc_4 == 16 : 
          (_th_blink_tid_324 == 5)? th_myfunc_5 == 16 : 
          (_th_blink_tid_324 == 6)? th_myfunc_6 == 16 : 
          (_th_blink_tid_324 == 7)? th_myfunc_7 == 16 : 
          (_th_blink_tid_324 == 8)? th_myfunc_8 == 16 : 
          (_th_blink_tid_324 == 9)? th_myfunc_9 == 16 : 
          (_th_blink_tid_324 == 10)? th_myfunc_10 == 16 : 
          (_th_blink_tid_324 == 11)? th_myfunc_11 == 16 : 
          (_th_blink_tid_324 == 12)? th_myfunc_12 == 16 : 
          (_th_blink_tid_324 == 13)? th_myfunc_13 == 16 : 
          (_th_blink_tid_324 == 14)? th_myfunc_14 == 16 : 
          (_th_blink_tid_324 == 15)? th_myfunc_15 == 16 : 
          (_th_blink_tid_324 == 16)? th_myfunc_16 == 16 : 
          (_th_blink_tid_324 == 17)? th_myfunc_17 == 16 : 
          (_th_blink_tid_324 == 18)? th_myfunc_18 == 16 : 
          (_th_blink_tid_324 == 19)? th_myfunc_19 == 16 : 
          (_th_blink_tid_324 == 20)? th_myfunc_20 == 16 : 
          (_th_blink_tid_324 == 21)? th_myfunc_21 == 16 : 
          (_th_blink_tid_324 == 22)? th_myfunc_22 == 16 : 
          (_th_blink_tid_324 == 23)? th_myfunc_23 == 16 : 
          (_th_blink_tid_324 == 24)? th_myfunc_24 == 16 : 
          (_th_blink_tid_324 == 25)? th_myfunc_25 == 16 : 
          (_th_blink_tid_324 == 26)? th_myfunc_26 == 16 : 
          (_th_blink_tid_324 == 27)? th_myfunc_27 == 16 : 
          (_th_blink_tid_324 == 28)? th_myfunc_28 == 16 : 
          (_th_blink_tid_324 == 29)? th_myfunc_29 == 16 : 
          (_th_blink_tid_324 == 30)? th_myfunc_30 == 16 : 
          (_th_blink_tid_324 == 31)? th_myfunc_31 == 16 : 
          (_th_blink_tid_324 == 32)? th_myfunc_32 == 16 : 
          (_th_blink_tid_324 == 33)? th_myfunc_33 == 16 : 
          (_th_blink_tid_324 == 34)? th_myfunc_34 == 16 : 
          (_th_blink_tid_324 == 35)? th_myfunc_35 == 16 : 
          (_th_blink_tid_324 == 36)? th_myfunc_36 == 16 : 
          (_th_blink_tid_324 == 37)? th_myfunc_37 == 16 : 
          (_th_blink_tid_324 == 38)? th_myfunc_38 == 16 : 
          (_th_blink_tid_324 == 39)? th_myfunc_39 == 16 : 
          (_th_blink_tid_324 == 40)? th_myfunc_40 == 16 : 
          (_th_blink_tid_324 == 41)? th_myfunc_41 == 16 : 
          (_th_blink_tid_324 == 42)? th_myfunc_42 == 16 : 
          (_th_blink_tid_324 == 43)? th_myfunc_43 == 16 : 
          (_th_blink_tid_324 == 44)? th_myfunc_44 == 16 : 
          (_th_blink_tid_324 == 45)? th_myfunc_45 == 16 : 
          (_th_blink_tid_324 == 46)? th_myfunc_46 == 16 : 
          (_th_blink_tid_324 == 47)? th_myfunc_47 == 16 : 
          (_th_blink_tid_324 == 48)? th_myfunc_48 == 16 : 
          (_th_blink_tid_324 == 49)? th_myfunc_49 == 16 : 
          (_th_blink_tid_324 == 50)? th_myfunc_50 == 16 : 
          (_th_blink_tid_324 == 51)? th_myfunc_51 == 16 : 
          (_th_blink_tid_324 == 52)? th_myfunc_52 == 16 : 
          (_th_blink_tid_324 == 53)? th_myfunc_53 == 16 : 
          (_th_blink_tid_324 == 54)? th_myfunc_54 == 16 : 
          (_th_blink_tid_324 == 55)? th_myfunc_55 == 16 : 
          (_th_blink_tid_324 == 56)? th_myfunc_56 == 16 : 
          (_th_blink_tid_324 == 57)? th_myfunc_57 == 16 : 
          (_th_blink_tid_324 == 58)? th_myfunc_58 == 16 : 
          (_th_blink_tid_324 == 59)? th_myfunc_59 == 16 : 
          (_th_blink_tid_324 == 60)? th_myfunc_60 == 16 : 
          (_th_blink_tid_324 == 61)? th_myfunc_61 == 16 : 
          (_th_blink_tid_324 == 62)? th_myfunc_62 == 16 : 
          (_th_blink_tid_324 == 63)? th_myfunc_63 == 16 : 0) begin
            th_blink <= th_blink_16;
          end 
        end
        th_blink_16: begin
          _th_blink_tid_324 <= _th_blink_tid_324 + 1;
          th_blink <= th_blink_14;
        end
        th_blink_17: begin
          _th_blink_tid_324 <= 0;
          th_blink <= th_blink_18;
        end
        th_blink_18: begin
          if(_th_blink_tid_324 < 64) begin
            th_blink <= th_blink_19;
          end else begin
            th_blink <= th_blink_20;
          end
        end
        th_blink_19: begin
          _th_blink_tid_324 <= _th_blink_tid_324 + 1;
          th_blink <= th_blink_18;
        end
        th_blink_20: begin
          done <= 1;
          th_blink <= th_blink_21;
        end
        th_blink_21: begin
          th_blink <= th_blink_2;
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count <= 0;
    end else begin
      if(th_blink == 1) begin
        count <= 0;
      end 
      if(th_myfunc_0 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_1 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_2 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_3 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_4 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_5 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_6 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_7 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_8 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_9 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_10 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_11 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_12 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_13 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_14 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_15 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_16 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_17 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_18 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_19 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_20 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_21 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_22 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_23 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_24 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_25 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_26 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_27 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_28 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_29 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_30 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_31 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_32 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_33 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_34 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_35 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_36 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_37 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_38 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_39 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_40 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_41 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_42 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_43 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_44 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_45 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_46 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_47 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_48 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_49 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_50 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_51 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_52 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_53 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_54 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_55 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_56 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_57 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_58 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_59 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_60 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_61 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_62 == 12) begin
        count <= count + 1;
      end 
      if(th_myfunc_63 == 12) begin
        count <= count + 1;
      end 
    end
  end

  localparam th_myfunc_0_1 = 1;
  localparam th_myfunc_0_2 = 2;
  localparam th_myfunc_0_3 = 3;
  localparam th_myfunc_0_4 = 4;
  localparam th_myfunc_0_5 = 5;
  localparam th_myfunc_0_6 = 6;
  localparam th_myfunc_0_7 = 7;
  localparam th_myfunc_0_8 = 8;
  localparam th_myfunc_0_9 = 9;
  localparam th_myfunc_0_10 = 10;
  localparam th_myfunc_0_11 = 11;
  localparam th_myfunc_0_12 = 12;
  localparam th_myfunc_0_13 = 13;
  localparam th_myfunc_0_14 = 14;
  localparam th_myfunc_0_15 = 15;
  localparam th_myfunc_0_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_0 <= th_myfunc_0_init;
      _th_myfunc_0_called <= 0;
      _th_myfunc_0_tid_325 <= 0;
      _th_myfunc_0_tid_326 <= 0;
      _th_myfunc_0_time_327 <= 0;
      _th_myfunc_0_i_328 <= 0;
      _th_myfunc_0___329 <= 0;
    end else begin
      case(th_myfunc_0)
        th_myfunc_0_init: begin
          if(_th_myfunc_start[0] && (th_blink == 10)) begin
            _th_myfunc_0_called <= 1;
          end 
          if(_th_myfunc_start[0] && (th_blink == 10)) begin
            _th_myfunc_0_tid_325 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[0]) begin
            th_myfunc_0 <= th_myfunc_0_1;
          end 
        end
        th_myfunc_0_1: begin
          _th_myfunc_0_tid_326 <= _th_myfunc_0_tid_325;
          th_myfunc_0 <= th_myfunc_0_2;
        end
        th_myfunc_0_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 0)) begin
            th_myfunc_0 <= th_myfunc_0_3;
          end 
        end
        th_myfunc_0_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 0))) begin
            th_myfunc_0 <= th_myfunc_0_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 0)) begin
            th_myfunc_0 <= th_myfunc_0_4;
          end 
        end
        th_myfunc_0_4: begin
          $display("Thread %d Lock", _th_myfunc_0_tid_326);
          th_myfunc_0 <= th_myfunc_0_5;
        end
        th_myfunc_0_5: begin
          _th_myfunc_0_time_327 <= sw;
          th_myfunc_0 <= th_myfunc_0_6;
        end
        th_myfunc_0_6: begin
          _th_myfunc_0_i_328 <= 0;
          th_myfunc_0 <= th_myfunc_0_7;
        end
        th_myfunc_0_7: begin
          if(_th_myfunc_0_i_328 < _th_myfunc_0_time_327) begin
            th_myfunc_0 <= th_myfunc_0_8;
          end else begin
            th_myfunc_0 <= th_myfunc_0_12;
          end
        end
        th_myfunc_0_8: begin
          _th_myfunc_0___329 <= 0;
          th_myfunc_0 <= th_myfunc_0_9;
        end
        th_myfunc_0_9: begin
          if(_th_myfunc_0___329 < 1024) begin
            th_myfunc_0 <= th_myfunc_0_10;
          end else begin
            th_myfunc_0 <= th_myfunc_0_11;
          end
        end
        th_myfunc_0_10: begin
          _th_myfunc_0___329 <= _th_myfunc_0___329 + 1;
          th_myfunc_0 <= th_myfunc_0_9;
        end
        th_myfunc_0_11: begin
          _th_myfunc_0_i_328 <= _th_myfunc_0_i_328 + 1;
          th_myfunc_0 <= th_myfunc_0_7;
        end
        th_myfunc_0_12: begin
          th_myfunc_0 <= th_myfunc_0_13;
        end
        th_myfunc_0_13: begin
          $display("Thread %d count = %d", _th_myfunc_0_tid_326, count);
          th_myfunc_0 <= th_myfunc_0_14;
        end
        th_myfunc_0_14: begin
          th_myfunc_0 <= th_myfunc_0_15;
        end
        th_myfunc_0_15: begin
          $display("Thread %d Unlock", _th_myfunc_0_tid_326);
          th_myfunc_0 <= th_myfunc_0_16;
        end
        th_myfunc_0_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 0)) begin
            _th_myfunc_0_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 0)) begin
            th_myfunc_0 <= th_myfunc_0_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_1_1 = 1;
  localparam th_myfunc_1_2 = 2;
  localparam th_myfunc_1_3 = 3;
  localparam th_myfunc_1_4 = 4;
  localparam th_myfunc_1_5 = 5;
  localparam th_myfunc_1_6 = 6;
  localparam th_myfunc_1_7 = 7;
  localparam th_myfunc_1_8 = 8;
  localparam th_myfunc_1_9 = 9;
  localparam th_myfunc_1_10 = 10;
  localparam th_myfunc_1_11 = 11;
  localparam th_myfunc_1_12 = 12;
  localparam th_myfunc_1_13 = 13;
  localparam th_myfunc_1_14 = 14;
  localparam th_myfunc_1_15 = 15;
  localparam th_myfunc_1_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_1 <= th_myfunc_1_init;
      _th_myfunc_1_called <= 0;
      _th_myfunc_1_tid_330 <= 0;
      _th_myfunc_1_tid_331 <= 0;
      _th_myfunc_1_time_332 <= 0;
      _th_myfunc_1_i_333 <= 0;
      _th_myfunc_1___334 <= 0;
    end else begin
      case(th_myfunc_1)
        th_myfunc_1_init: begin
          if(_th_myfunc_start[1] && (th_blink == 10)) begin
            _th_myfunc_1_called <= 1;
          end 
          if(_th_myfunc_start[1] && (th_blink == 10)) begin
            _th_myfunc_1_tid_330 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[1]) begin
            th_myfunc_1 <= th_myfunc_1_1;
          end 
        end
        th_myfunc_1_1: begin
          _th_myfunc_1_tid_331 <= _th_myfunc_1_tid_330;
          th_myfunc_1 <= th_myfunc_1_2;
        end
        th_myfunc_1_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 1)) begin
            th_myfunc_1 <= th_myfunc_1_3;
          end 
        end
        th_myfunc_1_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 1))) begin
            th_myfunc_1 <= th_myfunc_1_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 1)) begin
            th_myfunc_1 <= th_myfunc_1_4;
          end 
        end
        th_myfunc_1_4: begin
          $display("Thread %d Lock", _th_myfunc_1_tid_331);
          th_myfunc_1 <= th_myfunc_1_5;
        end
        th_myfunc_1_5: begin
          _th_myfunc_1_time_332 <= sw;
          th_myfunc_1 <= th_myfunc_1_6;
        end
        th_myfunc_1_6: begin
          _th_myfunc_1_i_333 <= 0;
          th_myfunc_1 <= th_myfunc_1_7;
        end
        th_myfunc_1_7: begin
          if(_th_myfunc_1_i_333 < _th_myfunc_1_time_332) begin
            th_myfunc_1 <= th_myfunc_1_8;
          end else begin
            th_myfunc_1 <= th_myfunc_1_12;
          end
        end
        th_myfunc_1_8: begin
          _th_myfunc_1___334 <= 0;
          th_myfunc_1 <= th_myfunc_1_9;
        end
        th_myfunc_1_9: begin
          if(_th_myfunc_1___334 < 1024) begin
            th_myfunc_1 <= th_myfunc_1_10;
          end else begin
            th_myfunc_1 <= th_myfunc_1_11;
          end
        end
        th_myfunc_1_10: begin
          _th_myfunc_1___334 <= _th_myfunc_1___334 + 1;
          th_myfunc_1 <= th_myfunc_1_9;
        end
        th_myfunc_1_11: begin
          _th_myfunc_1_i_333 <= _th_myfunc_1_i_333 + 1;
          th_myfunc_1 <= th_myfunc_1_7;
        end
        th_myfunc_1_12: begin
          th_myfunc_1 <= th_myfunc_1_13;
        end
        th_myfunc_1_13: begin
          $display("Thread %d count = %d", _th_myfunc_1_tid_331, count);
          th_myfunc_1 <= th_myfunc_1_14;
        end
        th_myfunc_1_14: begin
          th_myfunc_1 <= th_myfunc_1_15;
        end
        th_myfunc_1_15: begin
          $display("Thread %d Unlock", _th_myfunc_1_tid_331);
          th_myfunc_1 <= th_myfunc_1_16;
        end
        th_myfunc_1_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 1)) begin
            _th_myfunc_1_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 1)) begin
            th_myfunc_1 <= th_myfunc_1_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_2_1 = 1;
  localparam th_myfunc_2_2 = 2;
  localparam th_myfunc_2_3 = 3;
  localparam th_myfunc_2_4 = 4;
  localparam th_myfunc_2_5 = 5;
  localparam th_myfunc_2_6 = 6;
  localparam th_myfunc_2_7 = 7;
  localparam th_myfunc_2_8 = 8;
  localparam th_myfunc_2_9 = 9;
  localparam th_myfunc_2_10 = 10;
  localparam th_myfunc_2_11 = 11;
  localparam th_myfunc_2_12 = 12;
  localparam th_myfunc_2_13 = 13;
  localparam th_myfunc_2_14 = 14;
  localparam th_myfunc_2_15 = 15;
  localparam th_myfunc_2_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_2 <= th_myfunc_2_init;
      _th_myfunc_2_called <= 0;
      _th_myfunc_2_tid_335 <= 0;
      _th_myfunc_2_tid_336 <= 0;
      _th_myfunc_2_time_337 <= 0;
      _th_myfunc_2_i_338 <= 0;
      _th_myfunc_2___339 <= 0;
    end else begin
      case(th_myfunc_2)
        th_myfunc_2_init: begin
          if(_th_myfunc_start[2] && (th_blink == 10)) begin
            _th_myfunc_2_called <= 1;
          end 
          if(_th_myfunc_start[2] && (th_blink == 10)) begin
            _th_myfunc_2_tid_335 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[2]) begin
            th_myfunc_2 <= th_myfunc_2_1;
          end 
        end
        th_myfunc_2_1: begin
          _th_myfunc_2_tid_336 <= _th_myfunc_2_tid_335;
          th_myfunc_2 <= th_myfunc_2_2;
        end
        th_myfunc_2_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 2)) begin
            th_myfunc_2 <= th_myfunc_2_3;
          end 
        end
        th_myfunc_2_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 2))) begin
            th_myfunc_2 <= th_myfunc_2_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 2)) begin
            th_myfunc_2 <= th_myfunc_2_4;
          end 
        end
        th_myfunc_2_4: begin
          $display("Thread %d Lock", _th_myfunc_2_tid_336);
          th_myfunc_2 <= th_myfunc_2_5;
        end
        th_myfunc_2_5: begin
          _th_myfunc_2_time_337 <= sw;
          th_myfunc_2 <= th_myfunc_2_6;
        end
        th_myfunc_2_6: begin
          _th_myfunc_2_i_338 <= 0;
          th_myfunc_2 <= th_myfunc_2_7;
        end
        th_myfunc_2_7: begin
          if(_th_myfunc_2_i_338 < _th_myfunc_2_time_337) begin
            th_myfunc_2 <= th_myfunc_2_8;
          end else begin
            th_myfunc_2 <= th_myfunc_2_12;
          end
        end
        th_myfunc_2_8: begin
          _th_myfunc_2___339 <= 0;
          th_myfunc_2 <= th_myfunc_2_9;
        end
        th_myfunc_2_9: begin
          if(_th_myfunc_2___339 < 1024) begin
            th_myfunc_2 <= th_myfunc_2_10;
          end else begin
            th_myfunc_2 <= th_myfunc_2_11;
          end
        end
        th_myfunc_2_10: begin
          _th_myfunc_2___339 <= _th_myfunc_2___339 + 1;
          th_myfunc_2 <= th_myfunc_2_9;
        end
        th_myfunc_2_11: begin
          _th_myfunc_2_i_338 <= _th_myfunc_2_i_338 + 1;
          th_myfunc_2 <= th_myfunc_2_7;
        end
        th_myfunc_2_12: begin
          th_myfunc_2 <= th_myfunc_2_13;
        end
        th_myfunc_2_13: begin
          $display("Thread %d count = %d", _th_myfunc_2_tid_336, count);
          th_myfunc_2 <= th_myfunc_2_14;
        end
        th_myfunc_2_14: begin
          th_myfunc_2 <= th_myfunc_2_15;
        end
        th_myfunc_2_15: begin
          $display("Thread %d Unlock", _th_myfunc_2_tid_336);
          th_myfunc_2 <= th_myfunc_2_16;
        end
        th_myfunc_2_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 2)) begin
            _th_myfunc_2_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 2)) begin
            th_myfunc_2 <= th_myfunc_2_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_3_1 = 1;
  localparam th_myfunc_3_2 = 2;
  localparam th_myfunc_3_3 = 3;
  localparam th_myfunc_3_4 = 4;
  localparam th_myfunc_3_5 = 5;
  localparam th_myfunc_3_6 = 6;
  localparam th_myfunc_3_7 = 7;
  localparam th_myfunc_3_8 = 8;
  localparam th_myfunc_3_9 = 9;
  localparam th_myfunc_3_10 = 10;
  localparam th_myfunc_3_11 = 11;
  localparam th_myfunc_3_12 = 12;
  localparam th_myfunc_3_13 = 13;
  localparam th_myfunc_3_14 = 14;
  localparam th_myfunc_3_15 = 15;
  localparam th_myfunc_3_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_3 <= th_myfunc_3_init;
      _th_myfunc_3_called <= 0;
      _th_myfunc_3_tid_340 <= 0;
      _th_myfunc_3_tid_341 <= 0;
      _th_myfunc_3_time_342 <= 0;
      _th_myfunc_3_i_343 <= 0;
      _th_myfunc_3___344 <= 0;
    end else begin
      case(th_myfunc_3)
        th_myfunc_3_init: begin
          if(_th_myfunc_start[3] && (th_blink == 10)) begin
            _th_myfunc_3_called <= 1;
          end 
          if(_th_myfunc_start[3] && (th_blink == 10)) begin
            _th_myfunc_3_tid_340 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[3]) begin
            th_myfunc_3 <= th_myfunc_3_1;
          end 
        end
        th_myfunc_3_1: begin
          _th_myfunc_3_tid_341 <= _th_myfunc_3_tid_340;
          th_myfunc_3 <= th_myfunc_3_2;
        end
        th_myfunc_3_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 3)) begin
            th_myfunc_3 <= th_myfunc_3_3;
          end 
        end
        th_myfunc_3_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 3))) begin
            th_myfunc_3 <= th_myfunc_3_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 3)) begin
            th_myfunc_3 <= th_myfunc_3_4;
          end 
        end
        th_myfunc_3_4: begin
          $display("Thread %d Lock", _th_myfunc_3_tid_341);
          th_myfunc_3 <= th_myfunc_3_5;
        end
        th_myfunc_3_5: begin
          _th_myfunc_3_time_342 <= sw;
          th_myfunc_3 <= th_myfunc_3_6;
        end
        th_myfunc_3_6: begin
          _th_myfunc_3_i_343 <= 0;
          th_myfunc_3 <= th_myfunc_3_7;
        end
        th_myfunc_3_7: begin
          if(_th_myfunc_3_i_343 < _th_myfunc_3_time_342) begin
            th_myfunc_3 <= th_myfunc_3_8;
          end else begin
            th_myfunc_3 <= th_myfunc_3_12;
          end
        end
        th_myfunc_3_8: begin
          _th_myfunc_3___344 <= 0;
          th_myfunc_3 <= th_myfunc_3_9;
        end
        th_myfunc_3_9: begin
          if(_th_myfunc_3___344 < 1024) begin
            th_myfunc_3 <= th_myfunc_3_10;
          end else begin
            th_myfunc_3 <= th_myfunc_3_11;
          end
        end
        th_myfunc_3_10: begin
          _th_myfunc_3___344 <= _th_myfunc_3___344 + 1;
          th_myfunc_3 <= th_myfunc_3_9;
        end
        th_myfunc_3_11: begin
          _th_myfunc_3_i_343 <= _th_myfunc_3_i_343 + 1;
          th_myfunc_3 <= th_myfunc_3_7;
        end
        th_myfunc_3_12: begin
          th_myfunc_3 <= th_myfunc_3_13;
        end
        th_myfunc_3_13: begin
          $display("Thread %d count = %d", _th_myfunc_3_tid_341, count);
          th_myfunc_3 <= th_myfunc_3_14;
        end
        th_myfunc_3_14: begin
          th_myfunc_3 <= th_myfunc_3_15;
        end
        th_myfunc_3_15: begin
          $display("Thread %d Unlock", _th_myfunc_3_tid_341);
          th_myfunc_3 <= th_myfunc_3_16;
        end
        th_myfunc_3_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 3)) begin
            _th_myfunc_3_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 3)) begin
            th_myfunc_3 <= th_myfunc_3_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_4_1 = 1;
  localparam th_myfunc_4_2 = 2;
  localparam th_myfunc_4_3 = 3;
  localparam th_myfunc_4_4 = 4;
  localparam th_myfunc_4_5 = 5;
  localparam th_myfunc_4_6 = 6;
  localparam th_myfunc_4_7 = 7;
  localparam th_myfunc_4_8 = 8;
  localparam th_myfunc_4_9 = 9;
  localparam th_myfunc_4_10 = 10;
  localparam th_myfunc_4_11 = 11;
  localparam th_myfunc_4_12 = 12;
  localparam th_myfunc_4_13 = 13;
  localparam th_myfunc_4_14 = 14;
  localparam th_myfunc_4_15 = 15;
  localparam th_myfunc_4_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_4 <= th_myfunc_4_init;
      _th_myfunc_4_called <= 0;
      _th_myfunc_4_tid_345 <= 0;
      _th_myfunc_4_tid_346 <= 0;
      _th_myfunc_4_time_347 <= 0;
      _th_myfunc_4_i_348 <= 0;
      _th_myfunc_4___349 <= 0;
    end else begin
      case(th_myfunc_4)
        th_myfunc_4_init: begin
          if(_th_myfunc_start[4] && (th_blink == 10)) begin
            _th_myfunc_4_called <= 1;
          end 
          if(_th_myfunc_start[4] && (th_blink == 10)) begin
            _th_myfunc_4_tid_345 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[4]) begin
            th_myfunc_4 <= th_myfunc_4_1;
          end 
        end
        th_myfunc_4_1: begin
          _th_myfunc_4_tid_346 <= _th_myfunc_4_tid_345;
          th_myfunc_4 <= th_myfunc_4_2;
        end
        th_myfunc_4_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 4)) begin
            th_myfunc_4 <= th_myfunc_4_3;
          end 
        end
        th_myfunc_4_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 4))) begin
            th_myfunc_4 <= th_myfunc_4_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 4)) begin
            th_myfunc_4 <= th_myfunc_4_4;
          end 
        end
        th_myfunc_4_4: begin
          $display("Thread %d Lock", _th_myfunc_4_tid_346);
          th_myfunc_4 <= th_myfunc_4_5;
        end
        th_myfunc_4_5: begin
          _th_myfunc_4_time_347 <= sw;
          th_myfunc_4 <= th_myfunc_4_6;
        end
        th_myfunc_4_6: begin
          _th_myfunc_4_i_348 <= 0;
          th_myfunc_4 <= th_myfunc_4_7;
        end
        th_myfunc_4_7: begin
          if(_th_myfunc_4_i_348 < _th_myfunc_4_time_347) begin
            th_myfunc_4 <= th_myfunc_4_8;
          end else begin
            th_myfunc_4 <= th_myfunc_4_12;
          end
        end
        th_myfunc_4_8: begin
          _th_myfunc_4___349 <= 0;
          th_myfunc_4 <= th_myfunc_4_9;
        end
        th_myfunc_4_9: begin
          if(_th_myfunc_4___349 < 1024) begin
            th_myfunc_4 <= th_myfunc_4_10;
          end else begin
            th_myfunc_4 <= th_myfunc_4_11;
          end
        end
        th_myfunc_4_10: begin
          _th_myfunc_4___349 <= _th_myfunc_4___349 + 1;
          th_myfunc_4 <= th_myfunc_4_9;
        end
        th_myfunc_4_11: begin
          _th_myfunc_4_i_348 <= _th_myfunc_4_i_348 + 1;
          th_myfunc_4 <= th_myfunc_4_7;
        end
        th_myfunc_4_12: begin
          th_myfunc_4 <= th_myfunc_4_13;
        end
        th_myfunc_4_13: begin
          $display("Thread %d count = %d", _th_myfunc_4_tid_346, count);
          th_myfunc_4 <= th_myfunc_4_14;
        end
        th_myfunc_4_14: begin
          th_myfunc_4 <= th_myfunc_4_15;
        end
        th_myfunc_4_15: begin
          $display("Thread %d Unlock", _th_myfunc_4_tid_346);
          th_myfunc_4 <= th_myfunc_4_16;
        end
        th_myfunc_4_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 4)) begin
            _th_myfunc_4_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 4)) begin
            th_myfunc_4 <= th_myfunc_4_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_5_1 = 1;
  localparam th_myfunc_5_2 = 2;
  localparam th_myfunc_5_3 = 3;
  localparam th_myfunc_5_4 = 4;
  localparam th_myfunc_5_5 = 5;
  localparam th_myfunc_5_6 = 6;
  localparam th_myfunc_5_7 = 7;
  localparam th_myfunc_5_8 = 8;
  localparam th_myfunc_5_9 = 9;
  localparam th_myfunc_5_10 = 10;
  localparam th_myfunc_5_11 = 11;
  localparam th_myfunc_5_12 = 12;
  localparam th_myfunc_5_13 = 13;
  localparam th_myfunc_5_14 = 14;
  localparam th_myfunc_5_15 = 15;
  localparam th_myfunc_5_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_5 <= th_myfunc_5_init;
      _th_myfunc_5_called <= 0;
      _th_myfunc_5_tid_350 <= 0;
      _th_myfunc_5_tid_351 <= 0;
      _th_myfunc_5_time_352 <= 0;
      _th_myfunc_5_i_353 <= 0;
      _th_myfunc_5___354 <= 0;
    end else begin
      case(th_myfunc_5)
        th_myfunc_5_init: begin
          if(_th_myfunc_start[5] && (th_blink == 10)) begin
            _th_myfunc_5_called <= 1;
          end 
          if(_th_myfunc_start[5] && (th_blink == 10)) begin
            _th_myfunc_5_tid_350 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[5]) begin
            th_myfunc_5 <= th_myfunc_5_1;
          end 
        end
        th_myfunc_5_1: begin
          _th_myfunc_5_tid_351 <= _th_myfunc_5_tid_350;
          th_myfunc_5 <= th_myfunc_5_2;
        end
        th_myfunc_5_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 5)) begin
            th_myfunc_5 <= th_myfunc_5_3;
          end 
        end
        th_myfunc_5_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 5))) begin
            th_myfunc_5 <= th_myfunc_5_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 5)) begin
            th_myfunc_5 <= th_myfunc_5_4;
          end 
        end
        th_myfunc_5_4: begin
          $display("Thread %d Lock", _th_myfunc_5_tid_351);
          th_myfunc_5 <= th_myfunc_5_5;
        end
        th_myfunc_5_5: begin
          _th_myfunc_5_time_352 <= sw;
          th_myfunc_5 <= th_myfunc_5_6;
        end
        th_myfunc_5_6: begin
          _th_myfunc_5_i_353 <= 0;
          th_myfunc_5 <= th_myfunc_5_7;
        end
        th_myfunc_5_7: begin
          if(_th_myfunc_5_i_353 < _th_myfunc_5_time_352) begin
            th_myfunc_5 <= th_myfunc_5_8;
          end else begin
            th_myfunc_5 <= th_myfunc_5_12;
          end
        end
        th_myfunc_5_8: begin
          _th_myfunc_5___354 <= 0;
          th_myfunc_5 <= th_myfunc_5_9;
        end
        th_myfunc_5_9: begin
          if(_th_myfunc_5___354 < 1024) begin
            th_myfunc_5 <= th_myfunc_5_10;
          end else begin
            th_myfunc_5 <= th_myfunc_5_11;
          end
        end
        th_myfunc_5_10: begin
          _th_myfunc_5___354 <= _th_myfunc_5___354 + 1;
          th_myfunc_5 <= th_myfunc_5_9;
        end
        th_myfunc_5_11: begin
          _th_myfunc_5_i_353 <= _th_myfunc_5_i_353 + 1;
          th_myfunc_5 <= th_myfunc_5_7;
        end
        th_myfunc_5_12: begin
          th_myfunc_5 <= th_myfunc_5_13;
        end
        th_myfunc_5_13: begin
          $display("Thread %d count = %d", _th_myfunc_5_tid_351, count);
          th_myfunc_5 <= th_myfunc_5_14;
        end
        th_myfunc_5_14: begin
          th_myfunc_5 <= th_myfunc_5_15;
        end
        th_myfunc_5_15: begin
          $display("Thread %d Unlock", _th_myfunc_5_tid_351);
          th_myfunc_5 <= th_myfunc_5_16;
        end
        th_myfunc_5_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 5)) begin
            _th_myfunc_5_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 5)) begin
            th_myfunc_5 <= th_myfunc_5_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_6_1 = 1;
  localparam th_myfunc_6_2 = 2;
  localparam th_myfunc_6_3 = 3;
  localparam th_myfunc_6_4 = 4;
  localparam th_myfunc_6_5 = 5;
  localparam th_myfunc_6_6 = 6;
  localparam th_myfunc_6_7 = 7;
  localparam th_myfunc_6_8 = 8;
  localparam th_myfunc_6_9 = 9;
  localparam th_myfunc_6_10 = 10;
  localparam th_myfunc_6_11 = 11;
  localparam th_myfunc_6_12 = 12;
  localparam th_myfunc_6_13 = 13;
  localparam th_myfunc_6_14 = 14;
  localparam th_myfunc_6_15 = 15;
  localparam th_myfunc_6_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_6 <= th_myfunc_6_init;
      _th_myfunc_6_called <= 0;
      _th_myfunc_6_tid_355 <= 0;
      _th_myfunc_6_tid_356 <= 0;
      _th_myfunc_6_time_357 <= 0;
      _th_myfunc_6_i_358 <= 0;
      _th_myfunc_6___359 <= 0;
    end else begin
      case(th_myfunc_6)
        th_myfunc_6_init: begin
          if(_th_myfunc_start[6] && (th_blink == 10)) begin
            _th_myfunc_6_called <= 1;
          end 
          if(_th_myfunc_start[6] && (th_blink == 10)) begin
            _th_myfunc_6_tid_355 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[6]) begin
            th_myfunc_6 <= th_myfunc_6_1;
          end 
        end
        th_myfunc_6_1: begin
          _th_myfunc_6_tid_356 <= _th_myfunc_6_tid_355;
          th_myfunc_6 <= th_myfunc_6_2;
        end
        th_myfunc_6_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 6)) begin
            th_myfunc_6 <= th_myfunc_6_3;
          end 
        end
        th_myfunc_6_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 6))) begin
            th_myfunc_6 <= th_myfunc_6_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 6)) begin
            th_myfunc_6 <= th_myfunc_6_4;
          end 
        end
        th_myfunc_6_4: begin
          $display("Thread %d Lock", _th_myfunc_6_tid_356);
          th_myfunc_6 <= th_myfunc_6_5;
        end
        th_myfunc_6_5: begin
          _th_myfunc_6_time_357 <= sw;
          th_myfunc_6 <= th_myfunc_6_6;
        end
        th_myfunc_6_6: begin
          _th_myfunc_6_i_358 <= 0;
          th_myfunc_6 <= th_myfunc_6_7;
        end
        th_myfunc_6_7: begin
          if(_th_myfunc_6_i_358 < _th_myfunc_6_time_357) begin
            th_myfunc_6 <= th_myfunc_6_8;
          end else begin
            th_myfunc_6 <= th_myfunc_6_12;
          end
        end
        th_myfunc_6_8: begin
          _th_myfunc_6___359 <= 0;
          th_myfunc_6 <= th_myfunc_6_9;
        end
        th_myfunc_6_9: begin
          if(_th_myfunc_6___359 < 1024) begin
            th_myfunc_6 <= th_myfunc_6_10;
          end else begin
            th_myfunc_6 <= th_myfunc_6_11;
          end
        end
        th_myfunc_6_10: begin
          _th_myfunc_6___359 <= _th_myfunc_6___359 + 1;
          th_myfunc_6 <= th_myfunc_6_9;
        end
        th_myfunc_6_11: begin
          _th_myfunc_6_i_358 <= _th_myfunc_6_i_358 + 1;
          th_myfunc_6 <= th_myfunc_6_7;
        end
        th_myfunc_6_12: begin
          th_myfunc_6 <= th_myfunc_6_13;
        end
        th_myfunc_6_13: begin
          $display("Thread %d count = %d", _th_myfunc_6_tid_356, count);
          th_myfunc_6 <= th_myfunc_6_14;
        end
        th_myfunc_6_14: begin
          th_myfunc_6 <= th_myfunc_6_15;
        end
        th_myfunc_6_15: begin
          $display("Thread %d Unlock", _th_myfunc_6_tid_356);
          th_myfunc_6 <= th_myfunc_6_16;
        end
        th_myfunc_6_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 6)) begin
            _th_myfunc_6_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 6)) begin
            th_myfunc_6 <= th_myfunc_6_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_7_1 = 1;
  localparam th_myfunc_7_2 = 2;
  localparam th_myfunc_7_3 = 3;
  localparam th_myfunc_7_4 = 4;
  localparam th_myfunc_7_5 = 5;
  localparam th_myfunc_7_6 = 6;
  localparam th_myfunc_7_7 = 7;
  localparam th_myfunc_7_8 = 8;
  localparam th_myfunc_7_9 = 9;
  localparam th_myfunc_7_10 = 10;
  localparam th_myfunc_7_11 = 11;
  localparam th_myfunc_7_12 = 12;
  localparam th_myfunc_7_13 = 13;
  localparam th_myfunc_7_14 = 14;
  localparam th_myfunc_7_15 = 15;
  localparam th_myfunc_7_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_7 <= th_myfunc_7_init;
      _th_myfunc_7_called <= 0;
      _th_myfunc_7_tid_360 <= 0;
      _th_myfunc_7_tid_361 <= 0;
      _th_myfunc_7_time_362 <= 0;
      _th_myfunc_7_i_363 <= 0;
      _th_myfunc_7___364 <= 0;
    end else begin
      case(th_myfunc_7)
        th_myfunc_7_init: begin
          if(_th_myfunc_start[7] && (th_blink == 10)) begin
            _th_myfunc_7_called <= 1;
          end 
          if(_th_myfunc_start[7] && (th_blink == 10)) begin
            _th_myfunc_7_tid_360 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[7]) begin
            th_myfunc_7 <= th_myfunc_7_1;
          end 
        end
        th_myfunc_7_1: begin
          _th_myfunc_7_tid_361 <= _th_myfunc_7_tid_360;
          th_myfunc_7 <= th_myfunc_7_2;
        end
        th_myfunc_7_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 7)) begin
            th_myfunc_7 <= th_myfunc_7_3;
          end 
        end
        th_myfunc_7_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 7))) begin
            th_myfunc_7 <= th_myfunc_7_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 7)) begin
            th_myfunc_7 <= th_myfunc_7_4;
          end 
        end
        th_myfunc_7_4: begin
          $display("Thread %d Lock", _th_myfunc_7_tid_361);
          th_myfunc_7 <= th_myfunc_7_5;
        end
        th_myfunc_7_5: begin
          _th_myfunc_7_time_362 <= sw;
          th_myfunc_7 <= th_myfunc_7_6;
        end
        th_myfunc_7_6: begin
          _th_myfunc_7_i_363 <= 0;
          th_myfunc_7 <= th_myfunc_7_7;
        end
        th_myfunc_7_7: begin
          if(_th_myfunc_7_i_363 < _th_myfunc_7_time_362) begin
            th_myfunc_7 <= th_myfunc_7_8;
          end else begin
            th_myfunc_7 <= th_myfunc_7_12;
          end
        end
        th_myfunc_7_8: begin
          _th_myfunc_7___364 <= 0;
          th_myfunc_7 <= th_myfunc_7_9;
        end
        th_myfunc_7_9: begin
          if(_th_myfunc_7___364 < 1024) begin
            th_myfunc_7 <= th_myfunc_7_10;
          end else begin
            th_myfunc_7 <= th_myfunc_7_11;
          end
        end
        th_myfunc_7_10: begin
          _th_myfunc_7___364 <= _th_myfunc_7___364 + 1;
          th_myfunc_7 <= th_myfunc_7_9;
        end
        th_myfunc_7_11: begin
          _th_myfunc_7_i_363 <= _th_myfunc_7_i_363 + 1;
          th_myfunc_7 <= th_myfunc_7_7;
        end
        th_myfunc_7_12: begin
          th_myfunc_7 <= th_myfunc_7_13;
        end
        th_myfunc_7_13: begin
          $display("Thread %d count = %d", _th_myfunc_7_tid_361, count);
          th_myfunc_7 <= th_myfunc_7_14;
        end
        th_myfunc_7_14: begin
          th_myfunc_7 <= th_myfunc_7_15;
        end
        th_myfunc_7_15: begin
          $display("Thread %d Unlock", _th_myfunc_7_tid_361);
          th_myfunc_7 <= th_myfunc_7_16;
        end
        th_myfunc_7_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 7)) begin
            _th_myfunc_7_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 7)) begin
            th_myfunc_7 <= th_myfunc_7_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_8_1 = 1;
  localparam th_myfunc_8_2 = 2;
  localparam th_myfunc_8_3 = 3;
  localparam th_myfunc_8_4 = 4;
  localparam th_myfunc_8_5 = 5;
  localparam th_myfunc_8_6 = 6;
  localparam th_myfunc_8_7 = 7;
  localparam th_myfunc_8_8 = 8;
  localparam th_myfunc_8_9 = 9;
  localparam th_myfunc_8_10 = 10;
  localparam th_myfunc_8_11 = 11;
  localparam th_myfunc_8_12 = 12;
  localparam th_myfunc_8_13 = 13;
  localparam th_myfunc_8_14 = 14;
  localparam th_myfunc_8_15 = 15;
  localparam th_myfunc_8_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_8 <= th_myfunc_8_init;
      _th_myfunc_8_called <= 0;
      _th_myfunc_8_tid_365 <= 0;
      _th_myfunc_8_tid_366 <= 0;
      _th_myfunc_8_time_367 <= 0;
      _th_myfunc_8_i_368 <= 0;
      _th_myfunc_8___369 <= 0;
    end else begin
      case(th_myfunc_8)
        th_myfunc_8_init: begin
          if(_th_myfunc_start[8] && (th_blink == 10)) begin
            _th_myfunc_8_called <= 1;
          end 
          if(_th_myfunc_start[8] && (th_blink == 10)) begin
            _th_myfunc_8_tid_365 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[8]) begin
            th_myfunc_8 <= th_myfunc_8_1;
          end 
        end
        th_myfunc_8_1: begin
          _th_myfunc_8_tid_366 <= _th_myfunc_8_tid_365;
          th_myfunc_8 <= th_myfunc_8_2;
        end
        th_myfunc_8_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 8)) begin
            th_myfunc_8 <= th_myfunc_8_3;
          end 
        end
        th_myfunc_8_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 8))) begin
            th_myfunc_8 <= th_myfunc_8_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 8)) begin
            th_myfunc_8 <= th_myfunc_8_4;
          end 
        end
        th_myfunc_8_4: begin
          $display("Thread %d Lock", _th_myfunc_8_tid_366);
          th_myfunc_8 <= th_myfunc_8_5;
        end
        th_myfunc_8_5: begin
          _th_myfunc_8_time_367 <= sw;
          th_myfunc_8 <= th_myfunc_8_6;
        end
        th_myfunc_8_6: begin
          _th_myfunc_8_i_368 <= 0;
          th_myfunc_8 <= th_myfunc_8_7;
        end
        th_myfunc_8_7: begin
          if(_th_myfunc_8_i_368 < _th_myfunc_8_time_367) begin
            th_myfunc_8 <= th_myfunc_8_8;
          end else begin
            th_myfunc_8 <= th_myfunc_8_12;
          end
        end
        th_myfunc_8_8: begin
          _th_myfunc_8___369 <= 0;
          th_myfunc_8 <= th_myfunc_8_9;
        end
        th_myfunc_8_9: begin
          if(_th_myfunc_8___369 < 1024) begin
            th_myfunc_8 <= th_myfunc_8_10;
          end else begin
            th_myfunc_8 <= th_myfunc_8_11;
          end
        end
        th_myfunc_8_10: begin
          _th_myfunc_8___369 <= _th_myfunc_8___369 + 1;
          th_myfunc_8 <= th_myfunc_8_9;
        end
        th_myfunc_8_11: begin
          _th_myfunc_8_i_368 <= _th_myfunc_8_i_368 + 1;
          th_myfunc_8 <= th_myfunc_8_7;
        end
        th_myfunc_8_12: begin
          th_myfunc_8 <= th_myfunc_8_13;
        end
        th_myfunc_8_13: begin
          $display("Thread %d count = %d", _th_myfunc_8_tid_366, count);
          th_myfunc_8 <= th_myfunc_8_14;
        end
        th_myfunc_8_14: begin
          th_myfunc_8 <= th_myfunc_8_15;
        end
        th_myfunc_8_15: begin
          $display("Thread %d Unlock", _th_myfunc_8_tid_366);
          th_myfunc_8 <= th_myfunc_8_16;
        end
        th_myfunc_8_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 8)) begin
            _th_myfunc_8_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 8)) begin
            th_myfunc_8 <= th_myfunc_8_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_9_1 = 1;
  localparam th_myfunc_9_2 = 2;
  localparam th_myfunc_9_3 = 3;
  localparam th_myfunc_9_4 = 4;
  localparam th_myfunc_9_5 = 5;
  localparam th_myfunc_9_6 = 6;
  localparam th_myfunc_9_7 = 7;
  localparam th_myfunc_9_8 = 8;
  localparam th_myfunc_9_9 = 9;
  localparam th_myfunc_9_10 = 10;
  localparam th_myfunc_9_11 = 11;
  localparam th_myfunc_9_12 = 12;
  localparam th_myfunc_9_13 = 13;
  localparam th_myfunc_9_14 = 14;
  localparam th_myfunc_9_15 = 15;
  localparam th_myfunc_9_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_9 <= th_myfunc_9_init;
      _th_myfunc_9_called <= 0;
      _th_myfunc_9_tid_370 <= 0;
      _th_myfunc_9_tid_371 <= 0;
      _th_myfunc_9_time_372 <= 0;
      _th_myfunc_9_i_373 <= 0;
      _th_myfunc_9___374 <= 0;
    end else begin
      case(th_myfunc_9)
        th_myfunc_9_init: begin
          if(_th_myfunc_start[9] && (th_blink == 10)) begin
            _th_myfunc_9_called <= 1;
          end 
          if(_th_myfunc_start[9] && (th_blink == 10)) begin
            _th_myfunc_9_tid_370 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[9]) begin
            th_myfunc_9 <= th_myfunc_9_1;
          end 
        end
        th_myfunc_9_1: begin
          _th_myfunc_9_tid_371 <= _th_myfunc_9_tid_370;
          th_myfunc_9 <= th_myfunc_9_2;
        end
        th_myfunc_9_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 9)) begin
            th_myfunc_9 <= th_myfunc_9_3;
          end 
        end
        th_myfunc_9_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 9))) begin
            th_myfunc_9 <= th_myfunc_9_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 9)) begin
            th_myfunc_9 <= th_myfunc_9_4;
          end 
        end
        th_myfunc_9_4: begin
          $display("Thread %d Lock", _th_myfunc_9_tid_371);
          th_myfunc_9 <= th_myfunc_9_5;
        end
        th_myfunc_9_5: begin
          _th_myfunc_9_time_372 <= sw;
          th_myfunc_9 <= th_myfunc_9_6;
        end
        th_myfunc_9_6: begin
          _th_myfunc_9_i_373 <= 0;
          th_myfunc_9 <= th_myfunc_9_7;
        end
        th_myfunc_9_7: begin
          if(_th_myfunc_9_i_373 < _th_myfunc_9_time_372) begin
            th_myfunc_9 <= th_myfunc_9_8;
          end else begin
            th_myfunc_9 <= th_myfunc_9_12;
          end
        end
        th_myfunc_9_8: begin
          _th_myfunc_9___374 <= 0;
          th_myfunc_9 <= th_myfunc_9_9;
        end
        th_myfunc_9_9: begin
          if(_th_myfunc_9___374 < 1024) begin
            th_myfunc_9 <= th_myfunc_9_10;
          end else begin
            th_myfunc_9 <= th_myfunc_9_11;
          end
        end
        th_myfunc_9_10: begin
          _th_myfunc_9___374 <= _th_myfunc_9___374 + 1;
          th_myfunc_9 <= th_myfunc_9_9;
        end
        th_myfunc_9_11: begin
          _th_myfunc_9_i_373 <= _th_myfunc_9_i_373 + 1;
          th_myfunc_9 <= th_myfunc_9_7;
        end
        th_myfunc_9_12: begin
          th_myfunc_9 <= th_myfunc_9_13;
        end
        th_myfunc_9_13: begin
          $display("Thread %d count = %d", _th_myfunc_9_tid_371, count);
          th_myfunc_9 <= th_myfunc_9_14;
        end
        th_myfunc_9_14: begin
          th_myfunc_9 <= th_myfunc_9_15;
        end
        th_myfunc_9_15: begin
          $display("Thread %d Unlock", _th_myfunc_9_tid_371);
          th_myfunc_9 <= th_myfunc_9_16;
        end
        th_myfunc_9_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 9)) begin
            _th_myfunc_9_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 9)) begin
            th_myfunc_9 <= th_myfunc_9_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_10_1 = 1;
  localparam th_myfunc_10_2 = 2;
  localparam th_myfunc_10_3 = 3;
  localparam th_myfunc_10_4 = 4;
  localparam th_myfunc_10_5 = 5;
  localparam th_myfunc_10_6 = 6;
  localparam th_myfunc_10_7 = 7;
  localparam th_myfunc_10_8 = 8;
  localparam th_myfunc_10_9 = 9;
  localparam th_myfunc_10_10 = 10;
  localparam th_myfunc_10_11 = 11;
  localparam th_myfunc_10_12 = 12;
  localparam th_myfunc_10_13 = 13;
  localparam th_myfunc_10_14 = 14;
  localparam th_myfunc_10_15 = 15;
  localparam th_myfunc_10_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_10 <= th_myfunc_10_init;
      _th_myfunc_10_called <= 0;
      _th_myfunc_10_tid_375 <= 0;
      _th_myfunc_10_tid_376 <= 0;
      _th_myfunc_10_time_377 <= 0;
      _th_myfunc_10_i_378 <= 0;
      _th_myfunc_10___379 <= 0;
    end else begin
      case(th_myfunc_10)
        th_myfunc_10_init: begin
          if(_th_myfunc_start[10] && (th_blink == 10)) begin
            _th_myfunc_10_called <= 1;
          end 
          if(_th_myfunc_start[10] && (th_blink == 10)) begin
            _th_myfunc_10_tid_375 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[10]) begin
            th_myfunc_10 <= th_myfunc_10_1;
          end 
        end
        th_myfunc_10_1: begin
          _th_myfunc_10_tid_376 <= _th_myfunc_10_tid_375;
          th_myfunc_10 <= th_myfunc_10_2;
        end
        th_myfunc_10_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 10)) begin
            th_myfunc_10 <= th_myfunc_10_3;
          end 
        end
        th_myfunc_10_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 10))) begin
            th_myfunc_10 <= th_myfunc_10_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 10)) begin
            th_myfunc_10 <= th_myfunc_10_4;
          end 
        end
        th_myfunc_10_4: begin
          $display("Thread %d Lock", _th_myfunc_10_tid_376);
          th_myfunc_10 <= th_myfunc_10_5;
        end
        th_myfunc_10_5: begin
          _th_myfunc_10_time_377 <= sw;
          th_myfunc_10 <= th_myfunc_10_6;
        end
        th_myfunc_10_6: begin
          _th_myfunc_10_i_378 <= 0;
          th_myfunc_10 <= th_myfunc_10_7;
        end
        th_myfunc_10_7: begin
          if(_th_myfunc_10_i_378 < _th_myfunc_10_time_377) begin
            th_myfunc_10 <= th_myfunc_10_8;
          end else begin
            th_myfunc_10 <= th_myfunc_10_12;
          end
        end
        th_myfunc_10_8: begin
          _th_myfunc_10___379 <= 0;
          th_myfunc_10 <= th_myfunc_10_9;
        end
        th_myfunc_10_9: begin
          if(_th_myfunc_10___379 < 1024) begin
            th_myfunc_10 <= th_myfunc_10_10;
          end else begin
            th_myfunc_10 <= th_myfunc_10_11;
          end
        end
        th_myfunc_10_10: begin
          _th_myfunc_10___379 <= _th_myfunc_10___379 + 1;
          th_myfunc_10 <= th_myfunc_10_9;
        end
        th_myfunc_10_11: begin
          _th_myfunc_10_i_378 <= _th_myfunc_10_i_378 + 1;
          th_myfunc_10 <= th_myfunc_10_7;
        end
        th_myfunc_10_12: begin
          th_myfunc_10 <= th_myfunc_10_13;
        end
        th_myfunc_10_13: begin
          $display("Thread %d count = %d", _th_myfunc_10_tid_376, count);
          th_myfunc_10 <= th_myfunc_10_14;
        end
        th_myfunc_10_14: begin
          th_myfunc_10 <= th_myfunc_10_15;
        end
        th_myfunc_10_15: begin
          $display("Thread %d Unlock", _th_myfunc_10_tid_376);
          th_myfunc_10 <= th_myfunc_10_16;
        end
        th_myfunc_10_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 10)) begin
            _th_myfunc_10_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 10)) begin
            th_myfunc_10 <= th_myfunc_10_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_11_1 = 1;
  localparam th_myfunc_11_2 = 2;
  localparam th_myfunc_11_3 = 3;
  localparam th_myfunc_11_4 = 4;
  localparam th_myfunc_11_5 = 5;
  localparam th_myfunc_11_6 = 6;
  localparam th_myfunc_11_7 = 7;
  localparam th_myfunc_11_8 = 8;
  localparam th_myfunc_11_9 = 9;
  localparam th_myfunc_11_10 = 10;
  localparam th_myfunc_11_11 = 11;
  localparam th_myfunc_11_12 = 12;
  localparam th_myfunc_11_13 = 13;
  localparam th_myfunc_11_14 = 14;
  localparam th_myfunc_11_15 = 15;
  localparam th_myfunc_11_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_11 <= th_myfunc_11_init;
      _th_myfunc_11_called <= 0;
      _th_myfunc_11_tid_380 <= 0;
      _th_myfunc_11_tid_381 <= 0;
      _th_myfunc_11_time_382 <= 0;
      _th_myfunc_11_i_383 <= 0;
      _th_myfunc_11___384 <= 0;
    end else begin
      case(th_myfunc_11)
        th_myfunc_11_init: begin
          if(_th_myfunc_start[11] && (th_blink == 10)) begin
            _th_myfunc_11_called <= 1;
          end 
          if(_th_myfunc_start[11] && (th_blink == 10)) begin
            _th_myfunc_11_tid_380 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[11]) begin
            th_myfunc_11 <= th_myfunc_11_1;
          end 
        end
        th_myfunc_11_1: begin
          _th_myfunc_11_tid_381 <= _th_myfunc_11_tid_380;
          th_myfunc_11 <= th_myfunc_11_2;
        end
        th_myfunc_11_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 11)) begin
            th_myfunc_11 <= th_myfunc_11_3;
          end 
        end
        th_myfunc_11_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 11))) begin
            th_myfunc_11 <= th_myfunc_11_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 11)) begin
            th_myfunc_11 <= th_myfunc_11_4;
          end 
        end
        th_myfunc_11_4: begin
          $display("Thread %d Lock", _th_myfunc_11_tid_381);
          th_myfunc_11 <= th_myfunc_11_5;
        end
        th_myfunc_11_5: begin
          _th_myfunc_11_time_382 <= sw;
          th_myfunc_11 <= th_myfunc_11_6;
        end
        th_myfunc_11_6: begin
          _th_myfunc_11_i_383 <= 0;
          th_myfunc_11 <= th_myfunc_11_7;
        end
        th_myfunc_11_7: begin
          if(_th_myfunc_11_i_383 < _th_myfunc_11_time_382) begin
            th_myfunc_11 <= th_myfunc_11_8;
          end else begin
            th_myfunc_11 <= th_myfunc_11_12;
          end
        end
        th_myfunc_11_8: begin
          _th_myfunc_11___384 <= 0;
          th_myfunc_11 <= th_myfunc_11_9;
        end
        th_myfunc_11_9: begin
          if(_th_myfunc_11___384 < 1024) begin
            th_myfunc_11 <= th_myfunc_11_10;
          end else begin
            th_myfunc_11 <= th_myfunc_11_11;
          end
        end
        th_myfunc_11_10: begin
          _th_myfunc_11___384 <= _th_myfunc_11___384 + 1;
          th_myfunc_11 <= th_myfunc_11_9;
        end
        th_myfunc_11_11: begin
          _th_myfunc_11_i_383 <= _th_myfunc_11_i_383 + 1;
          th_myfunc_11 <= th_myfunc_11_7;
        end
        th_myfunc_11_12: begin
          th_myfunc_11 <= th_myfunc_11_13;
        end
        th_myfunc_11_13: begin
          $display("Thread %d count = %d", _th_myfunc_11_tid_381, count);
          th_myfunc_11 <= th_myfunc_11_14;
        end
        th_myfunc_11_14: begin
          th_myfunc_11 <= th_myfunc_11_15;
        end
        th_myfunc_11_15: begin
          $display("Thread %d Unlock", _th_myfunc_11_tid_381);
          th_myfunc_11 <= th_myfunc_11_16;
        end
        th_myfunc_11_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 11)) begin
            _th_myfunc_11_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 11)) begin
            th_myfunc_11 <= th_myfunc_11_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_12_1 = 1;
  localparam th_myfunc_12_2 = 2;
  localparam th_myfunc_12_3 = 3;
  localparam th_myfunc_12_4 = 4;
  localparam th_myfunc_12_5 = 5;
  localparam th_myfunc_12_6 = 6;
  localparam th_myfunc_12_7 = 7;
  localparam th_myfunc_12_8 = 8;
  localparam th_myfunc_12_9 = 9;
  localparam th_myfunc_12_10 = 10;
  localparam th_myfunc_12_11 = 11;
  localparam th_myfunc_12_12 = 12;
  localparam th_myfunc_12_13 = 13;
  localparam th_myfunc_12_14 = 14;
  localparam th_myfunc_12_15 = 15;
  localparam th_myfunc_12_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_12 <= th_myfunc_12_init;
      _th_myfunc_12_called <= 0;
      _th_myfunc_12_tid_385 <= 0;
      _th_myfunc_12_tid_386 <= 0;
      _th_myfunc_12_time_387 <= 0;
      _th_myfunc_12_i_388 <= 0;
      _th_myfunc_12___389 <= 0;
    end else begin
      case(th_myfunc_12)
        th_myfunc_12_init: begin
          if(_th_myfunc_start[12] && (th_blink == 10)) begin
            _th_myfunc_12_called <= 1;
          end 
          if(_th_myfunc_start[12] && (th_blink == 10)) begin
            _th_myfunc_12_tid_385 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[12]) begin
            th_myfunc_12 <= th_myfunc_12_1;
          end 
        end
        th_myfunc_12_1: begin
          _th_myfunc_12_tid_386 <= _th_myfunc_12_tid_385;
          th_myfunc_12 <= th_myfunc_12_2;
        end
        th_myfunc_12_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 12)) begin
            th_myfunc_12 <= th_myfunc_12_3;
          end 
        end
        th_myfunc_12_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 12))) begin
            th_myfunc_12 <= th_myfunc_12_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 12)) begin
            th_myfunc_12 <= th_myfunc_12_4;
          end 
        end
        th_myfunc_12_4: begin
          $display("Thread %d Lock", _th_myfunc_12_tid_386);
          th_myfunc_12 <= th_myfunc_12_5;
        end
        th_myfunc_12_5: begin
          _th_myfunc_12_time_387 <= sw;
          th_myfunc_12 <= th_myfunc_12_6;
        end
        th_myfunc_12_6: begin
          _th_myfunc_12_i_388 <= 0;
          th_myfunc_12 <= th_myfunc_12_7;
        end
        th_myfunc_12_7: begin
          if(_th_myfunc_12_i_388 < _th_myfunc_12_time_387) begin
            th_myfunc_12 <= th_myfunc_12_8;
          end else begin
            th_myfunc_12 <= th_myfunc_12_12;
          end
        end
        th_myfunc_12_8: begin
          _th_myfunc_12___389 <= 0;
          th_myfunc_12 <= th_myfunc_12_9;
        end
        th_myfunc_12_9: begin
          if(_th_myfunc_12___389 < 1024) begin
            th_myfunc_12 <= th_myfunc_12_10;
          end else begin
            th_myfunc_12 <= th_myfunc_12_11;
          end
        end
        th_myfunc_12_10: begin
          _th_myfunc_12___389 <= _th_myfunc_12___389 + 1;
          th_myfunc_12 <= th_myfunc_12_9;
        end
        th_myfunc_12_11: begin
          _th_myfunc_12_i_388 <= _th_myfunc_12_i_388 + 1;
          th_myfunc_12 <= th_myfunc_12_7;
        end
        th_myfunc_12_12: begin
          th_myfunc_12 <= th_myfunc_12_13;
        end
        th_myfunc_12_13: begin
          $display("Thread %d count = %d", _th_myfunc_12_tid_386, count);
          th_myfunc_12 <= th_myfunc_12_14;
        end
        th_myfunc_12_14: begin
          th_myfunc_12 <= th_myfunc_12_15;
        end
        th_myfunc_12_15: begin
          $display("Thread %d Unlock", _th_myfunc_12_tid_386);
          th_myfunc_12 <= th_myfunc_12_16;
        end
        th_myfunc_12_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 12)) begin
            _th_myfunc_12_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 12)) begin
            th_myfunc_12 <= th_myfunc_12_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_13_1 = 1;
  localparam th_myfunc_13_2 = 2;
  localparam th_myfunc_13_3 = 3;
  localparam th_myfunc_13_4 = 4;
  localparam th_myfunc_13_5 = 5;
  localparam th_myfunc_13_6 = 6;
  localparam th_myfunc_13_7 = 7;
  localparam th_myfunc_13_8 = 8;
  localparam th_myfunc_13_9 = 9;
  localparam th_myfunc_13_10 = 10;
  localparam th_myfunc_13_11 = 11;
  localparam th_myfunc_13_12 = 12;
  localparam th_myfunc_13_13 = 13;
  localparam th_myfunc_13_14 = 14;
  localparam th_myfunc_13_15 = 15;
  localparam th_myfunc_13_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_13 <= th_myfunc_13_init;
      _th_myfunc_13_called <= 0;
      _th_myfunc_13_tid_390 <= 0;
      _th_myfunc_13_tid_391 <= 0;
      _th_myfunc_13_time_392 <= 0;
      _th_myfunc_13_i_393 <= 0;
      _th_myfunc_13___394 <= 0;
    end else begin
      case(th_myfunc_13)
        th_myfunc_13_init: begin
          if(_th_myfunc_start[13] && (th_blink == 10)) begin
            _th_myfunc_13_called <= 1;
          end 
          if(_th_myfunc_start[13] && (th_blink == 10)) begin
            _th_myfunc_13_tid_390 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[13]) begin
            th_myfunc_13 <= th_myfunc_13_1;
          end 
        end
        th_myfunc_13_1: begin
          _th_myfunc_13_tid_391 <= _th_myfunc_13_tid_390;
          th_myfunc_13 <= th_myfunc_13_2;
        end
        th_myfunc_13_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 13)) begin
            th_myfunc_13 <= th_myfunc_13_3;
          end 
        end
        th_myfunc_13_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 13))) begin
            th_myfunc_13 <= th_myfunc_13_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 13)) begin
            th_myfunc_13 <= th_myfunc_13_4;
          end 
        end
        th_myfunc_13_4: begin
          $display("Thread %d Lock", _th_myfunc_13_tid_391);
          th_myfunc_13 <= th_myfunc_13_5;
        end
        th_myfunc_13_5: begin
          _th_myfunc_13_time_392 <= sw;
          th_myfunc_13 <= th_myfunc_13_6;
        end
        th_myfunc_13_6: begin
          _th_myfunc_13_i_393 <= 0;
          th_myfunc_13 <= th_myfunc_13_7;
        end
        th_myfunc_13_7: begin
          if(_th_myfunc_13_i_393 < _th_myfunc_13_time_392) begin
            th_myfunc_13 <= th_myfunc_13_8;
          end else begin
            th_myfunc_13 <= th_myfunc_13_12;
          end
        end
        th_myfunc_13_8: begin
          _th_myfunc_13___394 <= 0;
          th_myfunc_13 <= th_myfunc_13_9;
        end
        th_myfunc_13_9: begin
          if(_th_myfunc_13___394 < 1024) begin
            th_myfunc_13 <= th_myfunc_13_10;
          end else begin
            th_myfunc_13 <= th_myfunc_13_11;
          end
        end
        th_myfunc_13_10: begin
          _th_myfunc_13___394 <= _th_myfunc_13___394 + 1;
          th_myfunc_13 <= th_myfunc_13_9;
        end
        th_myfunc_13_11: begin
          _th_myfunc_13_i_393 <= _th_myfunc_13_i_393 + 1;
          th_myfunc_13 <= th_myfunc_13_7;
        end
        th_myfunc_13_12: begin
          th_myfunc_13 <= th_myfunc_13_13;
        end
        th_myfunc_13_13: begin
          $display("Thread %d count = %d", _th_myfunc_13_tid_391, count);
          th_myfunc_13 <= th_myfunc_13_14;
        end
        th_myfunc_13_14: begin
          th_myfunc_13 <= th_myfunc_13_15;
        end
        th_myfunc_13_15: begin
          $display("Thread %d Unlock", _th_myfunc_13_tid_391);
          th_myfunc_13 <= th_myfunc_13_16;
        end
        th_myfunc_13_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 13)) begin
            _th_myfunc_13_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 13)) begin
            th_myfunc_13 <= th_myfunc_13_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_14_1 = 1;
  localparam th_myfunc_14_2 = 2;
  localparam th_myfunc_14_3 = 3;
  localparam th_myfunc_14_4 = 4;
  localparam th_myfunc_14_5 = 5;
  localparam th_myfunc_14_6 = 6;
  localparam th_myfunc_14_7 = 7;
  localparam th_myfunc_14_8 = 8;
  localparam th_myfunc_14_9 = 9;
  localparam th_myfunc_14_10 = 10;
  localparam th_myfunc_14_11 = 11;
  localparam th_myfunc_14_12 = 12;
  localparam th_myfunc_14_13 = 13;
  localparam th_myfunc_14_14 = 14;
  localparam th_myfunc_14_15 = 15;
  localparam th_myfunc_14_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_14 <= th_myfunc_14_init;
      _th_myfunc_14_called <= 0;
      _th_myfunc_14_tid_395 <= 0;
      _th_myfunc_14_tid_396 <= 0;
      _th_myfunc_14_time_397 <= 0;
      _th_myfunc_14_i_398 <= 0;
      _th_myfunc_14___399 <= 0;
    end else begin
      case(th_myfunc_14)
        th_myfunc_14_init: begin
          if(_th_myfunc_start[14] && (th_blink == 10)) begin
            _th_myfunc_14_called <= 1;
          end 
          if(_th_myfunc_start[14] && (th_blink == 10)) begin
            _th_myfunc_14_tid_395 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[14]) begin
            th_myfunc_14 <= th_myfunc_14_1;
          end 
        end
        th_myfunc_14_1: begin
          _th_myfunc_14_tid_396 <= _th_myfunc_14_tid_395;
          th_myfunc_14 <= th_myfunc_14_2;
        end
        th_myfunc_14_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 14)) begin
            th_myfunc_14 <= th_myfunc_14_3;
          end 
        end
        th_myfunc_14_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 14))) begin
            th_myfunc_14 <= th_myfunc_14_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 14)) begin
            th_myfunc_14 <= th_myfunc_14_4;
          end 
        end
        th_myfunc_14_4: begin
          $display("Thread %d Lock", _th_myfunc_14_tid_396);
          th_myfunc_14 <= th_myfunc_14_5;
        end
        th_myfunc_14_5: begin
          _th_myfunc_14_time_397 <= sw;
          th_myfunc_14 <= th_myfunc_14_6;
        end
        th_myfunc_14_6: begin
          _th_myfunc_14_i_398 <= 0;
          th_myfunc_14 <= th_myfunc_14_7;
        end
        th_myfunc_14_7: begin
          if(_th_myfunc_14_i_398 < _th_myfunc_14_time_397) begin
            th_myfunc_14 <= th_myfunc_14_8;
          end else begin
            th_myfunc_14 <= th_myfunc_14_12;
          end
        end
        th_myfunc_14_8: begin
          _th_myfunc_14___399 <= 0;
          th_myfunc_14 <= th_myfunc_14_9;
        end
        th_myfunc_14_9: begin
          if(_th_myfunc_14___399 < 1024) begin
            th_myfunc_14 <= th_myfunc_14_10;
          end else begin
            th_myfunc_14 <= th_myfunc_14_11;
          end
        end
        th_myfunc_14_10: begin
          _th_myfunc_14___399 <= _th_myfunc_14___399 + 1;
          th_myfunc_14 <= th_myfunc_14_9;
        end
        th_myfunc_14_11: begin
          _th_myfunc_14_i_398 <= _th_myfunc_14_i_398 + 1;
          th_myfunc_14 <= th_myfunc_14_7;
        end
        th_myfunc_14_12: begin
          th_myfunc_14 <= th_myfunc_14_13;
        end
        th_myfunc_14_13: begin
          $display("Thread %d count = %d", _th_myfunc_14_tid_396, count);
          th_myfunc_14 <= th_myfunc_14_14;
        end
        th_myfunc_14_14: begin
          th_myfunc_14 <= th_myfunc_14_15;
        end
        th_myfunc_14_15: begin
          $display("Thread %d Unlock", _th_myfunc_14_tid_396);
          th_myfunc_14 <= th_myfunc_14_16;
        end
        th_myfunc_14_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 14)) begin
            _th_myfunc_14_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 14)) begin
            th_myfunc_14 <= th_myfunc_14_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_15_1 = 1;
  localparam th_myfunc_15_2 = 2;
  localparam th_myfunc_15_3 = 3;
  localparam th_myfunc_15_4 = 4;
  localparam th_myfunc_15_5 = 5;
  localparam th_myfunc_15_6 = 6;
  localparam th_myfunc_15_7 = 7;
  localparam th_myfunc_15_8 = 8;
  localparam th_myfunc_15_9 = 9;
  localparam th_myfunc_15_10 = 10;
  localparam th_myfunc_15_11 = 11;
  localparam th_myfunc_15_12 = 12;
  localparam th_myfunc_15_13 = 13;
  localparam th_myfunc_15_14 = 14;
  localparam th_myfunc_15_15 = 15;
  localparam th_myfunc_15_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_15 <= th_myfunc_15_init;
      _th_myfunc_15_called <= 0;
      _th_myfunc_15_tid_400 <= 0;
      _th_myfunc_15_tid_401 <= 0;
      _th_myfunc_15_time_402 <= 0;
      _th_myfunc_15_i_403 <= 0;
      _th_myfunc_15___404 <= 0;
    end else begin
      case(th_myfunc_15)
        th_myfunc_15_init: begin
          if(_th_myfunc_start[15] && (th_blink == 10)) begin
            _th_myfunc_15_called <= 1;
          end 
          if(_th_myfunc_start[15] && (th_blink == 10)) begin
            _th_myfunc_15_tid_400 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[15]) begin
            th_myfunc_15 <= th_myfunc_15_1;
          end 
        end
        th_myfunc_15_1: begin
          _th_myfunc_15_tid_401 <= _th_myfunc_15_tid_400;
          th_myfunc_15 <= th_myfunc_15_2;
        end
        th_myfunc_15_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 15)) begin
            th_myfunc_15 <= th_myfunc_15_3;
          end 
        end
        th_myfunc_15_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 15))) begin
            th_myfunc_15 <= th_myfunc_15_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 15)) begin
            th_myfunc_15 <= th_myfunc_15_4;
          end 
        end
        th_myfunc_15_4: begin
          $display("Thread %d Lock", _th_myfunc_15_tid_401);
          th_myfunc_15 <= th_myfunc_15_5;
        end
        th_myfunc_15_5: begin
          _th_myfunc_15_time_402 <= sw;
          th_myfunc_15 <= th_myfunc_15_6;
        end
        th_myfunc_15_6: begin
          _th_myfunc_15_i_403 <= 0;
          th_myfunc_15 <= th_myfunc_15_7;
        end
        th_myfunc_15_7: begin
          if(_th_myfunc_15_i_403 < _th_myfunc_15_time_402) begin
            th_myfunc_15 <= th_myfunc_15_8;
          end else begin
            th_myfunc_15 <= th_myfunc_15_12;
          end
        end
        th_myfunc_15_8: begin
          _th_myfunc_15___404 <= 0;
          th_myfunc_15 <= th_myfunc_15_9;
        end
        th_myfunc_15_9: begin
          if(_th_myfunc_15___404 < 1024) begin
            th_myfunc_15 <= th_myfunc_15_10;
          end else begin
            th_myfunc_15 <= th_myfunc_15_11;
          end
        end
        th_myfunc_15_10: begin
          _th_myfunc_15___404 <= _th_myfunc_15___404 + 1;
          th_myfunc_15 <= th_myfunc_15_9;
        end
        th_myfunc_15_11: begin
          _th_myfunc_15_i_403 <= _th_myfunc_15_i_403 + 1;
          th_myfunc_15 <= th_myfunc_15_7;
        end
        th_myfunc_15_12: begin
          th_myfunc_15 <= th_myfunc_15_13;
        end
        th_myfunc_15_13: begin
          $display("Thread %d count = %d", _th_myfunc_15_tid_401, count);
          th_myfunc_15 <= th_myfunc_15_14;
        end
        th_myfunc_15_14: begin
          th_myfunc_15 <= th_myfunc_15_15;
        end
        th_myfunc_15_15: begin
          $display("Thread %d Unlock", _th_myfunc_15_tid_401);
          th_myfunc_15 <= th_myfunc_15_16;
        end
        th_myfunc_15_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 15)) begin
            _th_myfunc_15_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 15)) begin
            th_myfunc_15 <= th_myfunc_15_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_16_1 = 1;
  localparam th_myfunc_16_2 = 2;
  localparam th_myfunc_16_3 = 3;
  localparam th_myfunc_16_4 = 4;
  localparam th_myfunc_16_5 = 5;
  localparam th_myfunc_16_6 = 6;
  localparam th_myfunc_16_7 = 7;
  localparam th_myfunc_16_8 = 8;
  localparam th_myfunc_16_9 = 9;
  localparam th_myfunc_16_10 = 10;
  localparam th_myfunc_16_11 = 11;
  localparam th_myfunc_16_12 = 12;
  localparam th_myfunc_16_13 = 13;
  localparam th_myfunc_16_14 = 14;
  localparam th_myfunc_16_15 = 15;
  localparam th_myfunc_16_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_16 <= th_myfunc_16_init;
      _th_myfunc_16_called <= 0;
      _th_myfunc_16_tid_405 <= 0;
      _th_myfunc_16_tid_406 <= 0;
      _th_myfunc_16_time_407 <= 0;
      _th_myfunc_16_i_408 <= 0;
      _th_myfunc_16___409 <= 0;
    end else begin
      case(th_myfunc_16)
        th_myfunc_16_init: begin
          if(_th_myfunc_start[16] && (th_blink == 10)) begin
            _th_myfunc_16_called <= 1;
          end 
          if(_th_myfunc_start[16] && (th_blink == 10)) begin
            _th_myfunc_16_tid_405 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[16]) begin
            th_myfunc_16 <= th_myfunc_16_1;
          end 
        end
        th_myfunc_16_1: begin
          _th_myfunc_16_tid_406 <= _th_myfunc_16_tid_405;
          th_myfunc_16 <= th_myfunc_16_2;
        end
        th_myfunc_16_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 16)) begin
            th_myfunc_16 <= th_myfunc_16_3;
          end 
        end
        th_myfunc_16_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 16))) begin
            th_myfunc_16 <= th_myfunc_16_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 16)) begin
            th_myfunc_16 <= th_myfunc_16_4;
          end 
        end
        th_myfunc_16_4: begin
          $display("Thread %d Lock", _th_myfunc_16_tid_406);
          th_myfunc_16 <= th_myfunc_16_5;
        end
        th_myfunc_16_5: begin
          _th_myfunc_16_time_407 <= sw;
          th_myfunc_16 <= th_myfunc_16_6;
        end
        th_myfunc_16_6: begin
          _th_myfunc_16_i_408 <= 0;
          th_myfunc_16 <= th_myfunc_16_7;
        end
        th_myfunc_16_7: begin
          if(_th_myfunc_16_i_408 < _th_myfunc_16_time_407) begin
            th_myfunc_16 <= th_myfunc_16_8;
          end else begin
            th_myfunc_16 <= th_myfunc_16_12;
          end
        end
        th_myfunc_16_8: begin
          _th_myfunc_16___409 <= 0;
          th_myfunc_16 <= th_myfunc_16_9;
        end
        th_myfunc_16_9: begin
          if(_th_myfunc_16___409 < 1024) begin
            th_myfunc_16 <= th_myfunc_16_10;
          end else begin
            th_myfunc_16 <= th_myfunc_16_11;
          end
        end
        th_myfunc_16_10: begin
          _th_myfunc_16___409 <= _th_myfunc_16___409 + 1;
          th_myfunc_16 <= th_myfunc_16_9;
        end
        th_myfunc_16_11: begin
          _th_myfunc_16_i_408 <= _th_myfunc_16_i_408 + 1;
          th_myfunc_16 <= th_myfunc_16_7;
        end
        th_myfunc_16_12: begin
          th_myfunc_16 <= th_myfunc_16_13;
        end
        th_myfunc_16_13: begin
          $display("Thread %d count = %d", _th_myfunc_16_tid_406, count);
          th_myfunc_16 <= th_myfunc_16_14;
        end
        th_myfunc_16_14: begin
          th_myfunc_16 <= th_myfunc_16_15;
        end
        th_myfunc_16_15: begin
          $display("Thread %d Unlock", _th_myfunc_16_tid_406);
          th_myfunc_16 <= th_myfunc_16_16;
        end
        th_myfunc_16_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 16)) begin
            _th_myfunc_16_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 16)) begin
            th_myfunc_16 <= th_myfunc_16_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_17_1 = 1;
  localparam th_myfunc_17_2 = 2;
  localparam th_myfunc_17_3 = 3;
  localparam th_myfunc_17_4 = 4;
  localparam th_myfunc_17_5 = 5;
  localparam th_myfunc_17_6 = 6;
  localparam th_myfunc_17_7 = 7;
  localparam th_myfunc_17_8 = 8;
  localparam th_myfunc_17_9 = 9;
  localparam th_myfunc_17_10 = 10;
  localparam th_myfunc_17_11 = 11;
  localparam th_myfunc_17_12 = 12;
  localparam th_myfunc_17_13 = 13;
  localparam th_myfunc_17_14 = 14;
  localparam th_myfunc_17_15 = 15;
  localparam th_myfunc_17_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_17 <= th_myfunc_17_init;
      _th_myfunc_17_called <= 0;
      _th_myfunc_17_tid_410 <= 0;
      _th_myfunc_17_tid_411 <= 0;
      _th_myfunc_17_time_412 <= 0;
      _th_myfunc_17_i_413 <= 0;
      _th_myfunc_17___414 <= 0;
    end else begin
      case(th_myfunc_17)
        th_myfunc_17_init: begin
          if(_th_myfunc_start[17] && (th_blink == 10)) begin
            _th_myfunc_17_called <= 1;
          end 
          if(_th_myfunc_start[17] && (th_blink == 10)) begin
            _th_myfunc_17_tid_410 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[17]) begin
            th_myfunc_17 <= th_myfunc_17_1;
          end 
        end
        th_myfunc_17_1: begin
          _th_myfunc_17_tid_411 <= _th_myfunc_17_tid_410;
          th_myfunc_17 <= th_myfunc_17_2;
        end
        th_myfunc_17_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 17)) begin
            th_myfunc_17 <= th_myfunc_17_3;
          end 
        end
        th_myfunc_17_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 17))) begin
            th_myfunc_17 <= th_myfunc_17_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 17)) begin
            th_myfunc_17 <= th_myfunc_17_4;
          end 
        end
        th_myfunc_17_4: begin
          $display("Thread %d Lock", _th_myfunc_17_tid_411);
          th_myfunc_17 <= th_myfunc_17_5;
        end
        th_myfunc_17_5: begin
          _th_myfunc_17_time_412 <= sw;
          th_myfunc_17 <= th_myfunc_17_6;
        end
        th_myfunc_17_6: begin
          _th_myfunc_17_i_413 <= 0;
          th_myfunc_17 <= th_myfunc_17_7;
        end
        th_myfunc_17_7: begin
          if(_th_myfunc_17_i_413 < _th_myfunc_17_time_412) begin
            th_myfunc_17 <= th_myfunc_17_8;
          end else begin
            th_myfunc_17 <= th_myfunc_17_12;
          end
        end
        th_myfunc_17_8: begin
          _th_myfunc_17___414 <= 0;
          th_myfunc_17 <= th_myfunc_17_9;
        end
        th_myfunc_17_9: begin
          if(_th_myfunc_17___414 < 1024) begin
            th_myfunc_17 <= th_myfunc_17_10;
          end else begin
            th_myfunc_17 <= th_myfunc_17_11;
          end
        end
        th_myfunc_17_10: begin
          _th_myfunc_17___414 <= _th_myfunc_17___414 + 1;
          th_myfunc_17 <= th_myfunc_17_9;
        end
        th_myfunc_17_11: begin
          _th_myfunc_17_i_413 <= _th_myfunc_17_i_413 + 1;
          th_myfunc_17 <= th_myfunc_17_7;
        end
        th_myfunc_17_12: begin
          th_myfunc_17 <= th_myfunc_17_13;
        end
        th_myfunc_17_13: begin
          $display("Thread %d count = %d", _th_myfunc_17_tid_411, count);
          th_myfunc_17 <= th_myfunc_17_14;
        end
        th_myfunc_17_14: begin
          th_myfunc_17 <= th_myfunc_17_15;
        end
        th_myfunc_17_15: begin
          $display("Thread %d Unlock", _th_myfunc_17_tid_411);
          th_myfunc_17 <= th_myfunc_17_16;
        end
        th_myfunc_17_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 17)) begin
            _th_myfunc_17_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 17)) begin
            th_myfunc_17 <= th_myfunc_17_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_18_1 = 1;
  localparam th_myfunc_18_2 = 2;
  localparam th_myfunc_18_3 = 3;
  localparam th_myfunc_18_4 = 4;
  localparam th_myfunc_18_5 = 5;
  localparam th_myfunc_18_6 = 6;
  localparam th_myfunc_18_7 = 7;
  localparam th_myfunc_18_8 = 8;
  localparam th_myfunc_18_9 = 9;
  localparam th_myfunc_18_10 = 10;
  localparam th_myfunc_18_11 = 11;
  localparam th_myfunc_18_12 = 12;
  localparam th_myfunc_18_13 = 13;
  localparam th_myfunc_18_14 = 14;
  localparam th_myfunc_18_15 = 15;
  localparam th_myfunc_18_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_18 <= th_myfunc_18_init;
      _th_myfunc_18_called <= 0;
      _th_myfunc_18_tid_415 <= 0;
      _th_myfunc_18_tid_416 <= 0;
      _th_myfunc_18_time_417 <= 0;
      _th_myfunc_18_i_418 <= 0;
      _th_myfunc_18___419 <= 0;
    end else begin
      case(th_myfunc_18)
        th_myfunc_18_init: begin
          if(_th_myfunc_start[18] && (th_blink == 10)) begin
            _th_myfunc_18_called <= 1;
          end 
          if(_th_myfunc_start[18] && (th_blink == 10)) begin
            _th_myfunc_18_tid_415 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[18]) begin
            th_myfunc_18 <= th_myfunc_18_1;
          end 
        end
        th_myfunc_18_1: begin
          _th_myfunc_18_tid_416 <= _th_myfunc_18_tid_415;
          th_myfunc_18 <= th_myfunc_18_2;
        end
        th_myfunc_18_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 18)) begin
            th_myfunc_18 <= th_myfunc_18_3;
          end 
        end
        th_myfunc_18_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 18))) begin
            th_myfunc_18 <= th_myfunc_18_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 18)) begin
            th_myfunc_18 <= th_myfunc_18_4;
          end 
        end
        th_myfunc_18_4: begin
          $display("Thread %d Lock", _th_myfunc_18_tid_416);
          th_myfunc_18 <= th_myfunc_18_5;
        end
        th_myfunc_18_5: begin
          _th_myfunc_18_time_417 <= sw;
          th_myfunc_18 <= th_myfunc_18_6;
        end
        th_myfunc_18_6: begin
          _th_myfunc_18_i_418 <= 0;
          th_myfunc_18 <= th_myfunc_18_7;
        end
        th_myfunc_18_7: begin
          if(_th_myfunc_18_i_418 < _th_myfunc_18_time_417) begin
            th_myfunc_18 <= th_myfunc_18_8;
          end else begin
            th_myfunc_18 <= th_myfunc_18_12;
          end
        end
        th_myfunc_18_8: begin
          _th_myfunc_18___419 <= 0;
          th_myfunc_18 <= th_myfunc_18_9;
        end
        th_myfunc_18_9: begin
          if(_th_myfunc_18___419 < 1024) begin
            th_myfunc_18 <= th_myfunc_18_10;
          end else begin
            th_myfunc_18 <= th_myfunc_18_11;
          end
        end
        th_myfunc_18_10: begin
          _th_myfunc_18___419 <= _th_myfunc_18___419 + 1;
          th_myfunc_18 <= th_myfunc_18_9;
        end
        th_myfunc_18_11: begin
          _th_myfunc_18_i_418 <= _th_myfunc_18_i_418 + 1;
          th_myfunc_18 <= th_myfunc_18_7;
        end
        th_myfunc_18_12: begin
          th_myfunc_18 <= th_myfunc_18_13;
        end
        th_myfunc_18_13: begin
          $display("Thread %d count = %d", _th_myfunc_18_tid_416, count);
          th_myfunc_18 <= th_myfunc_18_14;
        end
        th_myfunc_18_14: begin
          th_myfunc_18 <= th_myfunc_18_15;
        end
        th_myfunc_18_15: begin
          $display("Thread %d Unlock", _th_myfunc_18_tid_416);
          th_myfunc_18 <= th_myfunc_18_16;
        end
        th_myfunc_18_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 18)) begin
            _th_myfunc_18_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 18)) begin
            th_myfunc_18 <= th_myfunc_18_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_19_1 = 1;
  localparam th_myfunc_19_2 = 2;
  localparam th_myfunc_19_3 = 3;
  localparam th_myfunc_19_4 = 4;
  localparam th_myfunc_19_5 = 5;
  localparam th_myfunc_19_6 = 6;
  localparam th_myfunc_19_7 = 7;
  localparam th_myfunc_19_8 = 8;
  localparam th_myfunc_19_9 = 9;
  localparam th_myfunc_19_10 = 10;
  localparam th_myfunc_19_11 = 11;
  localparam th_myfunc_19_12 = 12;
  localparam th_myfunc_19_13 = 13;
  localparam th_myfunc_19_14 = 14;
  localparam th_myfunc_19_15 = 15;
  localparam th_myfunc_19_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_19 <= th_myfunc_19_init;
      _th_myfunc_19_called <= 0;
      _th_myfunc_19_tid_420 <= 0;
      _th_myfunc_19_tid_421 <= 0;
      _th_myfunc_19_time_422 <= 0;
      _th_myfunc_19_i_423 <= 0;
      _th_myfunc_19___424 <= 0;
    end else begin
      case(th_myfunc_19)
        th_myfunc_19_init: begin
          if(_th_myfunc_start[19] && (th_blink == 10)) begin
            _th_myfunc_19_called <= 1;
          end 
          if(_th_myfunc_start[19] && (th_blink == 10)) begin
            _th_myfunc_19_tid_420 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[19]) begin
            th_myfunc_19 <= th_myfunc_19_1;
          end 
        end
        th_myfunc_19_1: begin
          _th_myfunc_19_tid_421 <= _th_myfunc_19_tid_420;
          th_myfunc_19 <= th_myfunc_19_2;
        end
        th_myfunc_19_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 19)) begin
            th_myfunc_19 <= th_myfunc_19_3;
          end 
        end
        th_myfunc_19_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 19))) begin
            th_myfunc_19 <= th_myfunc_19_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 19)) begin
            th_myfunc_19 <= th_myfunc_19_4;
          end 
        end
        th_myfunc_19_4: begin
          $display("Thread %d Lock", _th_myfunc_19_tid_421);
          th_myfunc_19 <= th_myfunc_19_5;
        end
        th_myfunc_19_5: begin
          _th_myfunc_19_time_422 <= sw;
          th_myfunc_19 <= th_myfunc_19_6;
        end
        th_myfunc_19_6: begin
          _th_myfunc_19_i_423 <= 0;
          th_myfunc_19 <= th_myfunc_19_7;
        end
        th_myfunc_19_7: begin
          if(_th_myfunc_19_i_423 < _th_myfunc_19_time_422) begin
            th_myfunc_19 <= th_myfunc_19_8;
          end else begin
            th_myfunc_19 <= th_myfunc_19_12;
          end
        end
        th_myfunc_19_8: begin
          _th_myfunc_19___424 <= 0;
          th_myfunc_19 <= th_myfunc_19_9;
        end
        th_myfunc_19_9: begin
          if(_th_myfunc_19___424 < 1024) begin
            th_myfunc_19 <= th_myfunc_19_10;
          end else begin
            th_myfunc_19 <= th_myfunc_19_11;
          end
        end
        th_myfunc_19_10: begin
          _th_myfunc_19___424 <= _th_myfunc_19___424 + 1;
          th_myfunc_19 <= th_myfunc_19_9;
        end
        th_myfunc_19_11: begin
          _th_myfunc_19_i_423 <= _th_myfunc_19_i_423 + 1;
          th_myfunc_19 <= th_myfunc_19_7;
        end
        th_myfunc_19_12: begin
          th_myfunc_19 <= th_myfunc_19_13;
        end
        th_myfunc_19_13: begin
          $display("Thread %d count = %d", _th_myfunc_19_tid_421, count);
          th_myfunc_19 <= th_myfunc_19_14;
        end
        th_myfunc_19_14: begin
          th_myfunc_19 <= th_myfunc_19_15;
        end
        th_myfunc_19_15: begin
          $display("Thread %d Unlock", _th_myfunc_19_tid_421);
          th_myfunc_19 <= th_myfunc_19_16;
        end
        th_myfunc_19_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 19)) begin
            _th_myfunc_19_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 19)) begin
            th_myfunc_19 <= th_myfunc_19_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_20_1 = 1;
  localparam th_myfunc_20_2 = 2;
  localparam th_myfunc_20_3 = 3;
  localparam th_myfunc_20_4 = 4;
  localparam th_myfunc_20_5 = 5;
  localparam th_myfunc_20_6 = 6;
  localparam th_myfunc_20_7 = 7;
  localparam th_myfunc_20_8 = 8;
  localparam th_myfunc_20_9 = 9;
  localparam th_myfunc_20_10 = 10;
  localparam th_myfunc_20_11 = 11;
  localparam th_myfunc_20_12 = 12;
  localparam th_myfunc_20_13 = 13;
  localparam th_myfunc_20_14 = 14;
  localparam th_myfunc_20_15 = 15;
  localparam th_myfunc_20_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_20 <= th_myfunc_20_init;
      _th_myfunc_20_called <= 0;
      _th_myfunc_20_tid_425 <= 0;
      _th_myfunc_20_tid_426 <= 0;
      _th_myfunc_20_time_427 <= 0;
      _th_myfunc_20_i_428 <= 0;
      _th_myfunc_20___429 <= 0;
    end else begin
      case(th_myfunc_20)
        th_myfunc_20_init: begin
          if(_th_myfunc_start[20] && (th_blink == 10)) begin
            _th_myfunc_20_called <= 1;
          end 
          if(_th_myfunc_start[20] && (th_blink == 10)) begin
            _th_myfunc_20_tid_425 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[20]) begin
            th_myfunc_20 <= th_myfunc_20_1;
          end 
        end
        th_myfunc_20_1: begin
          _th_myfunc_20_tid_426 <= _th_myfunc_20_tid_425;
          th_myfunc_20 <= th_myfunc_20_2;
        end
        th_myfunc_20_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 20)) begin
            th_myfunc_20 <= th_myfunc_20_3;
          end 
        end
        th_myfunc_20_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 20))) begin
            th_myfunc_20 <= th_myfunc_20_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 20)) begin
            th_myfunc_20 <= th_myfunc_20_4;
          end 
        end
        th_myfunc_20_4: begin
          $display("Thread %d Lock", _th_myfunc_20_tid_426);
          th_myfunc_20 <= th_myfunc_20_5;
        end
        th_myfunc_20_5: begin
          _th_myfunc_20_time_427 <= sw;
          th_myfunc_20 <= th_myfunc_20_6;
        end
        th_myfunc_20_6: begin
          _th_myfunc_20_i_428 <= 0;
          th_myfunc_20 <= th_myfunc_20_7;
        end
        th_myfunc_20_7: begin
          if(_th_myfunc_20_i_428 < _th_myfunc_20_time_427) begin
            th_myfunc_20 <= th_myfunc_20_8;
          end else begin
            th_myfunc_20 <= th_myfunc_20_12;
          end
        end
        th_myfunc_20_8: begin
          _th_myfunc_20___429 <= 0;
          th_myfunc_20 <= th_myfunc_20_9;
        end
        th_myfunc_20_9: begin
          if(_th_myfunc_20___429 < 1024) begin
            th_myfunc_20 <= th_myfunc_20_10;
          end else begin
            th_myfunc_20 <= th_myfunc_20_11;
          end
        end
        th_myfunc_20_10: begin
          _th_myfunc_20___429 <= _th_myfunc_20___429 + 1;
          th_myfunc_20 <= th_myfunc_20_9;
        end
        th_myfunc_20_11: begin
          _th_myfunc_20_i_428 <= _th_myfunc_20_i_428 + 1;
          th_myfunc_20 <= th_myfunc_20_7;
        end
        th_myfunc_20_12: begin
          th_myfunc_20 <= th_myfunc_20_13;
        end
        th_myfunc_20_13: begin
          $display("Thread %d count = %d", _th_myfunc_20_tid_426, count);
          th_myfunc_20 <= th_myfunc_20_14;
        end
        th_myfunc_20_14: begin
          th_myfunc_20 <= th_myfunc_20_15;
        end
        th_myfunc_20_15: begin
          $display("Thread %d Unlock", _th_myfunc_20_tid_426);
          th_myfunc_20 <= th_myfunc_20_16;
        end
        th_myfunc_20_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 20)) begin
            _th_myfunc_20_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 20)) begin
            th_myfunc_20 <= th_myfunc_20_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_21_1 = 1;
  localparam th_myfunc_21_2 = 2;
  localparam th_myfunc_21_3 = 3;
  localparam th_myfunc_21_4 = 4;
  localparam th_myfunc_21_5 = 5;
  localparam th_myfunc_21_6 = 6;
  localparam th_myfunc_21_7 = 7;
  localparam th_myfunc_21_8 = 8;
  localparam th_myfunc_21_9 = 9;
  localparam th_myfunc_21_10 = 10;
  localparam th_myfunc_21_11 = 11;
  localparam th_myfunc_21_12 = 12;
  localparam th_myfunc_21_13 = 13;
  localparam th_myfunc_21_14 = 14;
  localparam th_myfunc_21_15 = 15;
  localparam th_myfunc_21_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_21 <= th_myfunc_21_init;
      _th_myfunc_21_called <= 0;
      _th_myfunc_21_tid_430 <= 0;
      _th_myfunc_21_tid_431 <= 0;
      _th_myfunc_21_time_432 <= 0;
      _th_myfunc_21_i_433 <= 0;
      _th_myfunc_21___434 <= 0;
    end else begin
      case(th_myfunc_21)
        th_myfunc_21_init: begin
          if(_th_myfunc_start[21] && (th_blink == 10)) begin
            _th_myfunc_21_called <= 1;
          end 
          if(_th_myfunc_start[21] && (th_blink == 10)) begin
            _th_myfunc_21_tid_430 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[21]) begin
            th_myfunc_21 <= th_myfunc_21_1;
          end 
        end
        th_myfunc_21_1: begin
          _th_myfunc_21_tid_431 <= _th_myfunc_21_tid_430;
          th_myfunc_21 <= th_myfunc_21_2;
        end
        th_myfunc_21_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 21)) begin
            th_myfunc_21 <= th_myfunc_21_3;
          end 
        end
        th_myfunc_21_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 21))) begin
            th_myfunc_21 <= th_myfunc_21_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 21)) begin
            th_myfunc_21 <= th_myfunc_21_4;
          end 
        end
        th_myfunc_21_4: begin
          $display("Thread %d Lock", _th_myfunc_21_tid_431);
          th_myfunc_21 <= th_myfunc_21_5;
        end
        th_myfunc_21_5: begin
          _th_myfunc_21_time_432 <= sw;
          th_myfunc_21 <= th_myfunc_21_6;
        end
        th_myfunc_21_6: begin
          _th_myfunc_21_i_433 <= 0;
          th_myfunc_21 <= th_myfunc_21_7;
        end
        th_myfunc_21_7: begin
          if(_th_myfunc_21_i_433 < _th_myfunc_21_time_432) begin
            th_myfunc_21 <= th_myfunc_21_8;
          end else begin
            th_myfunc_21 <= th_myfunc_21_12;
          end
        end
        th_myfunc_21_8: begin
          _th_myfunc_21___434 <= 0;
          th_myfunc_21 <= th_myfunc_21_9;
        end
        th_myfunc_21_9: begin
          if(_th_myfunc_21___434 < 1024) begin
            th_myfunc_21 <= th_myfunc_21_10;
          end else begin
            th_myfunc_21 <= th_myfunc_21_11;
          end
        end
        th_myfunc_21_10: begin
          _th_myfunc_21___434 <= _th_myfunc_21___434 + 1;
          th_myfunc_21 <= th_myfunc_21_9;
        end
        th_myfunc_21_11: begin
          _th_myfunc_21_i_433 <= _th_myfunc_21_i_433 + 1;
          th_myfunc_21 <= th_myfunc_21_7;
        end
        th_myfunc_21_12: begin
          th_myfunc_21 <= th_myfunc_21_13;
        end
        th_myfunc_21_13: begin
          $display("Thread %d count = %d", _th_myfunc_21_tid_431, count);
          th_myfunc_21 <= th_myfunc_21_14;
        end
        th_myfunc_21_14: begin
          th_myfunc_21 <= th_myfunc_21_15;
        end
        th_myfunc_21_15: begin
          $display("Thread %d Unlock", _th_myfunc_21_tid_431);
          th_myfunc_21 <= th_myfunc_21_16;
        end
        th_myfunc_21_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 21)) begin
            _th_myfunc_21_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 21)) begin
            th_myfunc_21 <= th_myfunc_21_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_22_1 = 1;
  localparam th_myfunc_22_2 = 2;
  localparam th_myfunc_22_3 = 3;
  localparam th_myfunc_22_4 = 4;
  localparam th_myfunc_22_5 = 5;
  localparam th_myfunc_22_6 = 6;
  localparam th_myfunc_22_7 = 7;
  localparam th_myfunc_22_8 = 8;
  localparam th_myfunc_22_9 = 9;
  localparam th_myfunc_22_10 = 10;
  localparam th_myfunc_22_11 = 11;
  localparam th_myfunc_22_12 = 12;
  localparam th_myfunc_22_13 = 13;
  localparam th_myfunc_22_14 = 14;
  localparam th_myfunc_22_15 = 15;
  localparam th_myfunc_22_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_22 <= th_myfunc_22_init;
      _th_myfunc_22_called <= 0;
      _th_myfunc_22_tid_435 <= 0;
      _th_myfunc_22_tid_436 <= 0;
      _th_myfunc_22_time_437 <= 0;
      _th_myfunc_22_i_438 <= 0;
      _th_myfunc_22___439 <= 0;
    end else begin
      case(th_myfunc_22)
        th_myfunc_22_init: begin
          if(_th_myfunc_start[22] && (th_blink == 10)) begin
            _th_myfunc_22_called <= 1;
          end 
          if(_th_myfunc_start[22] && (th_blink == 10)) begin
            _th_myfunc_22_tid_435 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[22]) begin
            th_myfunc_22 <= th_myfunc_22_1;
          end 
        end
        th_myfunc_22_1: begin
          _th_myfunc_22_tid_436 <= _th_myfunc_22_tid_435;
          th_myfunc_22 <= th_myfunc_22_2;
        end
        th_myfunc_22_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 22)) begin
            th_myfunc_22 <= th_myfunc_22_3;
          end 
        end
        th_myfunc_22_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 22))) begin
            th_myfunc_22 <= th_myfunc_22_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 22)) begin
            th_myfunc_22 <= th_myfunc_22_4;
          end 
        end
        th_myfunc_22_4: begin
          $display("Thread %d Lock", _th_myfunc_22_tid_436);
          th_myfunc_22 <= th_myfunc_22_5;
        end
        th_myfunc_22_5: begin
          _th_myfunc_22_time_437 <= sw;
          th_myfunc_22 <= th_myfunc_22_6;
        end
        th_myfunc_22_6: begin
          _th_myfunc_22_i_438 <= 0;
          th_myfunc_22 <= th_myfunc_22_7;
        end
        th_myfunc_22_7: begin
          if(_th_myfunc_22_i_438 < _th_myfunc_22_time_437) begin
            th_myfunc_22 <= th_myfunc_22_8;
          end else begin
            th_myfunc_22 <= th_myfunc_22_12;
          end
        end
        th_myfunc_22_8: begin
          _th_myfunc_22___439 <= 0;
          th_myfunc_22 <= th_myfunc_22_9;
        end
        th_myfunc_22_9: begin
          if(_th_myfunc_22___439 < 1024) begin
            th_myfunc_22 <= th_myfunc_22_10;
          end else begin
            th_myfunc_22 <= th_myfunc_22_11;
          end
        end
        th_myfunc_22_10: begin
          _th_myfunc_22___439 <= _th_myfunc_22___439 + 1;
          th_myfunc_22 <= th_myfunc_22_9;
        end
        th_myfunc_22_11: begin
          _th_myfunc_22_i_438 <= _th_myfunc_22_i_438 + 1;
          th_myfunc_22 <= th_myfunc_22_7;
        end
        th_myfunc_22_12: begin
          th_myfunc_22 <= th_myfunc_22_13;
        end
        th_myfunc_22_13: begin
          $display("Thread %d count = %d", _th_myfunc_22_tid_436, count);
          th_myfunc_22 <= th_myfunc_22_14;
        end
        th_myfunc_22_14: begin
          th_myfunc_22 <= th_myfunc_22_15;
        end
        th_myfunc_22_15: begin
          $display("Thread %d Unlock", _th_myfunc_22_tid_436);
          th_myfunc_22 <= th_myfunc_22_16;
        end
        th_myfunc_22_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 22)) begin
            _th_myfunc_22_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 22)) begin
            th_myfunc_22 <= th_myfunc_22_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_23_1 = 1;
  localparam th_myfunc_23_2 = 2;
  localparam th_myfunc_23_3 = 3;
  localparam th_myfunc_23_4 = 4;
  localparam th_myfunc_23_5 = 5;
  localparam th_myfunc_23_6 = 6;
  localparam th_myfunc_23_7 = 7;
  localparam th_myfunc_23_8 = 8;
  localparam th_myfunc_23_9 = 9;
  localparam th_myfunc_23_10 = 10;
  localparam th_myfunc_23_11 = 11;
  localparam th_myfunc_23_12 = 12;
  localparam th_myfunc_23_13 = 13;
  localparam th_myfunc_23_14 = 14;
  localparam th_myfunc_23_15 = 15;
  localparam th_myfunc_23_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_23 <= th_myfunc_23_init;
      _th_myfunc_23_called <= 0;
      _th_myfunc_23_tid_440 <= 0;
      _th_myfunc_23_tid_441 <= 0;
      _th_myfunc_23_time_442 <= 0;
      _th_myfunc_23_i_443 <= 0;
      _th_myfunc_23___444 <= 0;
    end else begin
      case(th_myfunc_23)
        th_myfunc_23_init: begin
          if(_th_myfunc_start[23] && (th_blink == 10)) begin
            _th_myfunc_23_called <= 1;
          end 
          if(_th_myfunc_start[23] && (th_blink == 10)) begin
            _th_myfunc_23_tid_440 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[23]) begin
            th_myfunc_23 <= th_myfunc_23_1;
          end 
        end
        th_myfunc_23_1: begin
          _th_myfunc_23_tid_441 <= _th_myfunc_23_tid_440;
          th_myfunc_23 <= th_myfunc_23_2;
        end
        th_myfunc_23_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 23)) begin
            th_myfunc_23 <= th_myfunc_23_3;
          end 
        end
        th_myfunc_23_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 23))) begin
            th_myfunc_23 <= th_myfunc_23_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 23)) begin
            th_myfunc_23 <= th_myfunc_23_4;
          end 
        end
        th_myfunc_23_4: begin
          $display("Thread %d Lock", _th_myfunc_23_tid_441);
          th_myfunc_23 <= th_myfunc_23_5;
        end
        th_myfunc_23_5: begin
          _th_myfunc_23_time_442 <= sw;
          th_myfunc_23 <= th_myfunc_23_6;
        end
        th_myfunc_23_6: begin
          _th_myfunc_23_i_443 <= 0;
          th_myfunc_23 <= th_myfunc_23_7;
        end
        th_myfunc_23_7: begin
          if(_th_myfunc_23_i_443 < _th_myfunc_23_time_442) begin
            th_myfunc_23 <= th_myfunc_23_8;
          end else begin
            th_myfunc_23 <= th_myfunc_23_12;
          end
        end
        th_myfunc_23_8: begin
          _th_myfunc_23___444 <= 0;
          th_myfunc_23 <= th_myfunc_23_9;
        end
        th_myfunc_23_9: begin
          if(_th_myfunc_23___444 < 1024) begin
            th_myfunc_23 <= th_myfunc_23_10;
          end else begin
            th_myfunc_23 <= th_myfunc_23_11;
          end
        end
        th_myfunc_23_10: begin
          _th_myfunc_23___444 <= _th_myfunc_23___444 + 1;
          th_myfunc_23 <= th_myfunc_23_9;
        end
        th_myfunc_23_11: begin
          _th_myfunc_23_i_443 <= _th_myfunc_23_i_443 + 1;
          th_myfunc_23 <= th_myfunc_23_7;
        end
        th_myfunc_23_12: begin
          th_myfunc_23 <= th_myfunc_23_13;
        end
        th_myfunc_23_13: begin
          $display("Thread %d count = %d", _th_myfunc_23_tid_441, count);
          th_myfunc_23 <= th_myfunc_23_14;
        end
        th_myfunc_23_14: begin
          th_myfunc_23 <= th_myfunc_23_15;
        end
        th_myfunc_23_15: begin
          $display("Thread %d Unlock", _th_myfunc_23_tid_441);
          th_myfunc_23 <= th_myfunc_23_16;
        end
        th_myfunc_23_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 23)) begin
            _th_myfunc_23_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 23)) begin
            th_myfunc_23 <= th_myfunc_23_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_24_1 = 1;
  localparam th_myfunc_24_2 = 2;
  localparam th_myfunc_24_3 = 3;
  localparam th_myfunc_24_4 = 4;
  localparam th_myfunc_24_5 = 5;
  localparam th_myfunc_24_6 = 6;
  localparam th_myfunc_24_7 = 7;
  localparam th_myfunc_24_8 = 8;
  localparam th_myfunc_24_9 = 9;
  localparam th_myfunc_24_10 = 10;
  localparam th_myfunc_24_11 = 11;
  localparam th_myfunc_24_12 = 12;
  localparam th_myfunc_24_13 = 13;
  localparam th_myfunc_24_14 = 14;
  localparam th_myfunc_24_15 = 15;
  localparam th_myfunc_24_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_24 <= th_myfunc_24_init;
      _th_myfunc_24_called <= 0;
      _th_myfunc_24_tid_445 <= 0;
      _th_myfunc_24_tid_446 <= 0;
      _th_myfunc_24_time_447 <= 0;
      _th_myfunc_24_i_448 <= 0;
      _th_myfunc_24___449 <= 0;
    end else begin
      case(th_myfunc_24)
        th_myfunc_24_init: begin
          if(_th_myfunc_start[24] && (th_blink == 10)) begin
            _th_myfunc_24_called <= 1;
          end 
          if(_th_myfunc_start[24] && (th_blink == 10)) begin
            _th_myfunc_24_tid_445 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[24]) begin
            th_myfunc_24 <= th_myfunc_24_1;
          end 
        end
        th_myfunc_24_1: begin
          _th_myfunc_24_tid_446 <= _th_myfunc_24_tid_445;
          th_myfunc_24 <= th_myfunc_24_2;
        end
        th_myfunc_24_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 24)) begin
            th_myfunc_24 <= th_myfunc_24_3;
          end 
        end
        th_myfunc_24_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 24))) begin
            th_myfunc_24 <= th_myfunc_24_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 24)) begin
            th_myfunc_24 <= th_myfunc_24_4;
          end 
        end
        th_myfunc_24_4: begin
          $display("Thread %d Lock", _th_myfunc_24_tid_446);
          th_myfunc_24 <= th_myfunc_24_5;
        end
        th_myfunc_24_5: begin
          _th_myfunc_24_time_447 <= sw;
          th_myfunc_24 <= th_myfunc_24_6;
        end
        th_myfunc_24_6: begin
          _th_myfunc_24_i_448 <= 0;
          th_myfunc_24 <= th_myfunc_24_7;
        end
        th_myfunc_24_7: begin
          if(_th_myfunc_24_i_448 < _th_myfunc_24_time_447) begin
            th_myfunc_24 <= th_myfunc_24_8;
          end else begin
            th_myfunc_24 <= th_myfunc_24_12;
          end
        end
        th_myfunc_24_8: begin
          _th_myfunc_24___449 <= 0;
          th_myfunc_24 <= th_myfunc_24_9;
        end
        th_myfunc_24_9: begin
          if(_th_myfunc_24___449 < 1024) begin
            th_myfunc_24 <= th_myfunc_24_10;
          end else begin
            th_myfunc_24 <= th_myfunc_24_11;
          end
        end
        th_myfunc_24_10: begin
          _th_myfunc_24___449 <= _th_myfunc_24___449 + 1;
          th_myfunc_24 <= th_myfunc_24_9;
        end
        th_myfunc_24_11: begin
          _th_myfunc_24_i_448 <= _th_myfunc_24_i_448 + 1;
          th_myfunc_24 <= th_myfunc_24_7;
        end
        th_myfunc_24_12: begin
          th_myfunc_24 <= th_myfunc_24_13;
        end
        th_myfunc_24_13: begin
          $display("Thread %d count = %d", _th_myfunc_24_tid_446, count);
          th_myfunc_24 <= th_myfunc_24_14;
        end
        th_myfunc_24_14: begin
          th_myfunc_24 <= th_myfunc_24_15;
        end
        th_myfunc_24_15: begin
          $display("Thread %d Unlock", _th_myfunc_24_tid_446);
          th_myfunc_24 <= th_myfunc_24_16;
        end
        th_myfunc_24_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 24)) begin
            _th_myfunc_24_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 24)) begin
            th_myfunc_24 <= th_myfunc_24_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_25_1 = 1;
  localparam th_myfunc_25_2 = 2;
  localparam th_myfunc_25_3 = 3;
  localparam th_myfunc_25_4 = 4;
  localparam th_myfunc_25_5 = 5;
  localparam th_myfunc_25_6 = 6;
  localparam th_myfunc_25_7 = 7;
  localparam th_myfunc_25_8 = 8;
  localparam th_myfunc_25_9 = 9;
  localparam th_myfunc_25_10 = 10;
  localparam th_myfunc_25_11 = 11;
  localparam th_myfunc_25_12 = 12;
  localparam th_myfunc_25_13 = 13;
  localparam th_myfunc_25_14 = 14;
  localparam th_myfunc_25_15 = 15;
  localparam th_myfunc_25_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_25 <= th_myfunc_25_init;
      _th_myfunc_25_called <= 0;
      _th_myfunc_25_tid_450 <= 0;
      _th_myfunc_25_tid_451 <= 0;
      _th_myfunc_25_time_452 <= 0;
      _th_myfunc_25_i_453 <= 0;
      _th_myfunc_25___454 <= 0;
    end else begin
      case(th_myfunc_25)
        th_myfunc_25_init: begin
          if(_th_myfunc_start[25] && (th_blink == 10)) begin
            _th_myfunc_25_called <= 1;
          end 
          if(_th_myfunc_start[25] && (th_blink == 10)) begin
            _th_myfunc_25_tid_450 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[25]) begin
            th_myfunc_25 <= th_myfunc_25_1;
          end 
        end
        th_myfunc_25_1: begin
          _th_myfunc_25_tid_451 <= _th_myfunc_25_tid_450;
          th_myfunc_25 <= th_myfunc_25_2;
        end
        th_myfunc_25_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 25)) begin
            th_myfunc_25 <= th_myfunc_25_3;
          end 
        end
        th_myfunc_25_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 25))) begin
            th_myfunc_25 <= th_myfunc_25_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 25)) begin
            th_myfunc_25 <= th_myfunc_25_4;
          end 
        end
        th_myfunc_25_4: begin
          $display("Thread %d Lock", _th_myfunc_25_tid_451);
          th_myfunc_25 <= th_myfunc_25_5;
        end
        th_myfunc_25_5: begin
          _th_myfunc_25_time_452 <= sw;
          th_myfunc_25 <= th_myfunc_25_6;
        end
        th_myfunc_25_6: begin
          _th_myfunc_25_i_453 <= 0;
          th_myfunc_25 <= th_myfunc_25_7;
        end
        th_myfunc_25_7: begin
          if(_th_myfunc_25_i_453 < _th_myfunc_25_time_452) begin
            th_myfunc_25 <= th_myfunc_25_8;
          end else begin
            th_myfunc_25 <= th_myfunc_25_12;
          end
        end
        th_myfunc_25_8: begin
          _th_myfunc_25___454 <= 0;
          th_myfunc_25 <= th_myfunc_25_9;
        end
        th_myfunc_25_9: begin
          if(_th_myfunc_25___454 < 1024) begin
            th_myfunc_25 <= th_myfunc_25_10;
          end else begin
            th_myfunc_25 <= th_myfunc_25_11;
          end
        end
        th_myfunc_25_10: begin
          _th_myfunc_25___454 <= _th_myfunc_25___454 + 1;
          th_myfunc_25 <= th_myfunc_25_9;
        end
        th_myfunc_25_11: begin
          _th_myfunc_25_i_453 <= _th_myfunc_25_i_453 + 1;
          th_myfunc_25 <= th_myfunc_25_7;
        end
        th_myfunc_25_12: begin
          th_myfunc_25 <= th_myfunc_25_13;
        end
        th_myfunc_25_13: begin
          $display("Thread %d count = %d", _th_myfunc_25_tid_451, count);
          th_myfunc_25 <= th_myfunc_25_14;
        end
        th_myfunc_25_14: begin
          th_myfunc_25 <= th_myfunc_25_15;
        end
        th_myfunc_25_15: begin
          $display("Thread %d Unlock", _th_myfunc_25_tid_451);
          th_myfunc_25 <= th_myfunc_25_16;
        end
        th_myfunc_25_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 25)) begin
            _th_myfunc_25_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 25)) begin
            th_myfunc_25 <= th_myfunc_25_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_26_1 = 1;
  localparam th_myfunc_26_2 = 2;
  localparam th_myfunc_26_3 = 3;
  localparam th_myfunc_26_4 = 4;
  localparam th_myfunc_26_5 = 5;
  localparam th_myfunc_26_6 = 6;
  localparam th_myfunc_26_7 = 7;
  localparam th_myfunc_26_8 = 8;
  localparam th_myfunc_26_9 = 9;
  localparam th_myfunc_26_10 = 10;
  localparam th_myfunc_26_11 = 11;
  localparam th_myfunc_26_12 = 12;
  localparam th_myfunc_26_13 = 13;
  localparam th_myfunc_26_14 = 14;
  localparam th_myfunc_26_15 = 15;
  localparam th_myfunc_26_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_26 <= th_myfunc_26_init;
      _th_myfunc_26_called <= 0;
      _th_myfunc_26_tid_455 <= 0;
      _th_myfunc_26_tid_456 <= 0;
      _th_myfunc_26_time_457 <= 0;
      _th_myfunc_26_i_458 <= 0;
      _th_myfunc_26___459 <= 0;
    end else begin
      case(th_myfunc_26)
        th_myfunc_26_init: begin
          if(_th_myfunc_start[26] && (th_blink == 10)) begin
            _th_myfunc_26_called <= 1;
          end 
          if(_th_myfunc_start[26] && (th_blink == 10)) begin
            _th_myfunc_26_tid_455 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[26]) begin
            th_myfunc_26 <= th_myfunc_26_1;
          end 
        end
        th_myfunc_26_1: begin
          _th_myfunc_26_tid_456 <= _th_myfunc_26_tid_455;
          th_myfunc_26 <= th_myfunc_26_2;
        end
        th_myfunc_26_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 26)) begin
            th_myfunc_26 <= th_myfunc_26_3;
          end 
        end
        th_myfunc_26_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 26))) begin
            th_myfunc_26 <= th_myfunc_26_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 26)) begin
            th_myfunc_26 <= th_myfunc_26_4;
          end 
        end
        th_myfunc_26_4: begin
          $display("Thread %d Lock", _th_myfunc_26_tid_456);
          th_myfunc_26 <= th_myfunc_26_5;
        end
        th_myfunc_26_5: begin
          _th_myfunc_26_time_457 <= sw;
          th_myfunc_26 <= th_myfunc_26_6;
        end
        th_myfunc_26_6: begin
          _th_myfunc_26_i_458 <= 0;
          th_myfunc_26 <= th_myfunc_26_7;
        end
        th_myfunc_26_7: begin
          if(_th_myfunc_26_i_458 < _th_myfunc_26_time_457) begin
            th_myfunc_26 <= th_myfunc_26_8;
          end else begin
            th_myfunc_26 <= th_myfunc_26_12;
          end
        end
        th_myfunc_26_8: begin
          _th_myfunc_26___459 <= 0;
          th_myfunc_26 <= th_myfunc_26_9;
        end
        th_myfunc_26_9: begin
          if(_th_myfunc_26___459 < 1024) begin
            th_myfunc_26 <= th_myfunc_26_10;
          end else begin
            th_myfunc_26 <= th_myfunc_26_11;
          end
        end
        th_myfunc_26_10: begin
          _th_myfunc_26___459 <= _th_myfunc_26___459 + 1;
          th_myfunc_26 <= th_myfunc_26_9;
        end
        th_myfunc_26_11: begin
          _th_myfunc_26_i_458 <= _th_myfunc_26_i_458 + 1;
          th_myfunc_26 <= th_myfunc_26_7;
        end
        th_myfunc_26_12: begin
          th_myfunc_26 <= th_myfunc_26_13;
        end
        th_myfunc_26_13: begin
          $display("Thread %d count = %d", _th_myfunc_26_tid_456, count);
          th_myfunc_26 <= th_myfunc_26_14;
        end
        th_myfunc_26_14: begin
          th_myfunc_26 <= th_myfunc_26_15;
        end
        th_myfunc_26_15: begin
          $display("Thread %d Unlock", _th_myfunc_26_tid_456);
          th_myfunc_26 <= th_myfunc_26_16;
        end
        th_myfunc_26_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 26)) begin
            _th_myfunc_26_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 26)) begin
            th_myfunc_26 <= th_myfunc_26_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_27_1 = 1;
  localparam th_myfunc_27_2 = 2;
  localparam th_myfunc_27_3 = 3;
  localparam th_myfunc_27_4 = 4;
  localparam th_myfunc_27_5 = 5;
  localparam th_myfunc_27_6 = 6;
  localparam th_myfunc_27_7 = 7;
  localparam th_myfunc_27_8 = 8;
  localparam th_myfunc_27_9 = 9;
  localparam th_myfunc_27_10 = 10;
  localparam th_myfunc_27_11 = 11;
  localparam th_myfunc_27_12 = 12;
  localparam th_myfunc_27_13 = 13;
  localparam th_myfunc_27_14 = 14;
  localparam th_myfunc_27_15 = 15;
  localparam th_myfunc_27_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_27 <= th_myfunc_27_init;
      _th_myfunc_27_called <= 0;
      _th_myfunc_27_tid_460 <= 0;
      _th_myfunc_27_tid_461 <= 0;
      _th_myfunc_27_time_462 <= 0;
      _th_myfunc_27_i_463 <= 0;
      _th_myfunc_27___464 <= 0;
    end else begin
      case(th_myfunc_27)
        th_myfunc_27_init: begin
          if(_th_myfunc_start[27] && (th_blink == 10)) begin
            _th_myfunc_27_called <= 1;
          end 
          if(_th_myfunc_start[27] && (th_blink == 10)) begin
            _th_myfunc_27_tid_460 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[27]) begin
            th_myfunc_27 <= th_myfunc_27_1;
          end 
        end
        th_myfunc_27_1: begin
          _th_myfunc_27_tid_461 <= _th_myfunc_27_tid_460;
          th_myfunc_27 <= th_myfunc_27_2;
        end
        th_myfunc_27_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 27)) begin
            th_myfunc_27 <= th_myfunc_27_3;
          end 
        end
        th_myfunc_27_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 27))) begin
            th_myfunc_27 <= th_myfunc_27_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 27)) begin
            th_myfunc_27 <= th_myfunc_27_4;
          end 
        end
        th_myfunc_27_4: begin
          $display("Thread %d Lock", _th_myfunc_27_tid_461);
          th_myfunc_27 <= th_myfunc_27_5;
        end
        th_myfunc_27_5: begin
          _th_myfunc_27_time_462 <= sw;
          th_myfunc_27 <= th_myfunc_27_6;
        end
        th_myfunc_27_6: begin
          _th_myfunc_27_i_463 <= 0;
          th_myfunc_27 <= th_myfunc_27_7;
        end
        th_myfunc_27_7: begin
          if(_th_myfunc_27_i_463 < _th_myfunc_27_time_462) begin
            th_myfunc_27 <= th_myfunc_27_8;
          end else begin
            th_myfunc_27 <= th_myfunc_27_12;
          end
        end
        th_myfunc_27_8: begin
          _th_myfunc_27___464 <= 0;
          th_myfunc_27 <= th_myfunc_27_9;
        end
        th_myfunc_27_9: begin
          if(_th_myfunc_27___464 < 1024) begin
            th_myfunc_27 <= th_myfunc_27_10;
          end else begin
            th_myfunc_27 <= th_myfunc_27_11;
          end
        end
        th_myfunc_27_10: begin
          _th_myfunc_27___464 <= _th_myfunc_27___464 + 1;
          th_myfunc_27 <= th_myfunc_27_9;
        end
        th_myfunc_27_11: begin
          _th_myfunc_27_i_463 <= _th_myfunc_27_i_463 + 1;
          th_myfunc_27 <= th_myfunc_27_7;
        end
        th_myfunc_27_12: begin
          th_myfunc_27 <= th_myfunc_27_13;
        end
        th_myfunc_27_13: begin
          $display("Thread %d count = %d", _th_myfunc_27_tid_461, count);
          th_myfunc_27 <= th_myfunc_27_14;
        end
        th_myfunc_27_14: begin
          th_myfunc_27 <= th_myfunc_27_15;
        end
        th_myfunc_27_15: begin
          $display("Thread %d Unlock", _th_myfunc_27_tid_461);
          th_myfunc_27 <= th_myfunc_27_16;
        end
        th_myfunc_27_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 27)) begin
            _th_myfunc_27_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 27)) begin
            th_myfunc_27 <= th_myfunc_27_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_28_1 = 1;
  localparam th_myfunc_28_2 = 2;
  localparam th_myfunc_28_3 = 3;
  localparam th_myfunc_28_4 = 4;
  localparam th_myfunc_28_5 = 5;
  localparam th_myfunc_28_6 = 6;
  localparam th_myfunc_28_7 = 7;
  localparam th_myfunc_28_8 = 8;
  localparam th_myfunc_28_9 = 9;
  localparam th_myfunc_28_10 = 10;
  localparam th_myfunc_28_11 = 11;
  localparam th_myfunc_28_12 = 12;
  localparam th_myfunc_28_13 = 13;
  localparam th_myfunc_28_14 = 14;
  localparam th_myfunc_28_15 = 15;
  localparam th_myfunc_28_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_28 <= th_myfunc_28_init;
      _th_myfunc_28_called <= 0;
      _th_myfunc_28_tid_465 <= 0;
      _th_myfunc_28_tid_466 <= 0;
      _th_myfunc_28_time_467 <= 0;
      _th_myfunc_28_i_468 <= 0;
      _th_myfunc_28___469 <= 0;
    end else begin
      case(th_myfunc_28)
        th_myfunc_28_init: begin
          if(_th_myfunc_start[28] && (th_blink == 10)) begin
            _th_myfunc_28_called <= 1;
          end 
          if(_th_myfunc_start[28] && (th_blink == 10)) begin
            _th_myfunc_28_tid_465 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[28]) begin
            th_myfunc_28 <= th_myfunc_28_1;
          end 
        end
        th_myfunc_28_1: begin
          _th_myfunc_28_tid_466 <= _th_myfunc_28_tid_465;
          th_myfunc_28 <= th_myfunc_28_2;
        end
        th_myfunc_28_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 28)) begin
            th_myfunc_28 <= th_myfunc_28_3;
          end 
        end
        th_myfunc_28_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 28))) begin
            th_myfunc_28 <= th_myfunc_28_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 28)) begin
            th_myfunc_28 <= th_myfunc_28_4;
          end 
        end
        th_myfunc_28_4: begin
          $display("Thread %d Lock", _th_myfunc_28_tid_466);
          th_myfunc_28 <= th_myfunc_28_5;
        end
        th_myfunc_28_5: begin
          _th_myfunc_28_time_467 <= sw;
          th_myfunc_28 <= th_myfunc_28_6;
        end
        th_myfunc_28_6: begin
          _th_myfunc_28_i_468 <= 0;
          th_myfunc_28 <= th_myfunc_28_7;
        end
        th_myfunc_28_7: begin
          if(_th_myfunc_28_i_468 < _th_myfunc_28_time_467) begin
            th_myfunc_28 <= th_myfunc_28_8;
          end else begin
            th_myfunc_28 <= th_myfunc_28_12;
          end
        end
        th_myfunc_28_8: begin
          _th_myfunc_28___469 <= 0;
          th_myfunc_28 <= th_myfunc_28_9;
        end
        th_myfunc_28_9: begin
          if(_th_myfunc_28___469 < 1024) begin
            th_myfunc_28 <= th_myfunc_28_10;
          end else begin
            th_myfunc_28 <= th_myfunc_28_11;
          end
        end
        th_myfunc_28_10: begin
          _th_myfunc_28___469 <= _th_myfunc_28___469 + 1;
          th_myfunc_28 <= th_myfunc_28_9;
        end
        th_myfunc_28_11: begin
          _th_myfunc_28_i_468 <= _th_myfunc_28_i_468 + 1;
          th_myfunc_28 <= th_myfunc_28_7;
        end
        th_myfunc_28_12: begin
          th_myfunc_28 <= th_myfunc_28_13;
        end
        th_myfunc_28_13: begin
          $display("Thread %d count = %d", _th_myfunc_28_tid_466, count);
          th_myfunc_28 <= th_myfunc_28_14;
        end
        th_myfunc_28_14: begin
          th_myfunc_28 <= th_myfunc_28_15;
        end
        th_myfunc_28_15: begin
          $display("Thread %d Unlock", _th_myfunc_28_tid_466);
          th_myfunc_28 <= th_myfunc_28_16;
        end
        th_myfunc_28_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 28)) begin
            _th_myfunc_28_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 28)) begin
            th_myfunc_28 <= th_myfunc_28_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_29_1 = 1;
  localparam th_myfunc_29_2 = 2;
  localparam th_myfunc_29_3 = 3;
  localparam th_myfunc_29_4 = 4;
  localparam th_myfunc_29_5 = 5;
  localparam th_myfunc_29_6 = 6;
  localparam th_myfunc_29_7 = 7;
  localparam th_myfunc_29_8 = 8;
  localparam th_myfunc_29_9 = 9;
  localparam th_myfunc_29_10 = 10;
  localparam th_myfunc_29_11 = 11;
  localparam th_myfunc_29_12 = 12;
  localparam th_myfunc_29_13 = 13;
  localparam th_myfunc_29_14 = 14;
  localparam th_myfunc_29_15 = 15;
  localparam th_myfunc_29_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_29 <= th_myfunc_29_init;
      _th_myfunc_29_called <= 0;
      _th_myfunc_29_tid_470 <= 0;
      _th_myfunc_29_tid_471 <= 0;
      _th_myfunc_29_time_472 <= 0;
      _th_myfunc_29_i_473 <= 0;
      _th_myfunc_29___474 <= 0;
    end else begin
      case(th_myfunc_29)
        th_myfunc_29_init: begin
          if(_th_myfunc_start[29] && (th_blink == 10)) begin
            _th_myfunc_29_called <= 1;
          end 
          if(_th_myfunc_start[29] && (th_blink == 10)) begin
            _th_myfunc_29_tid_470 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[29]) begin
            th_myfunc_29 <= th_myfunc_29_1;
          end 
        end
        th_myfunc_29_1: begin
          _th_myfunc_29_tid_471 <= _th_myfunc_29_tid_470;
          th_myfunc_29 <= th_myfunc_29_2;
        end
        th_myfunc_29_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 29)) begin
            th_myfunc_29 <= th_myfunc_29_3;
          end 
        end
        th_myfunc_29_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 29))) begin
            th_myfunc_29 <= th_myfunc_29_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 29)) begin
            th_myfunc_29 <= th_myfunc_29_4;
          end 
        end
        th_myfunc_29_4: begin
          $display("Thread %d Lock", _th_myfunc_29_tid_471);
          th_myfunc_29 <= th_myfunc_29_5;
        end
        th_myfunc_29_5: begin
          _th_myfunc_29_time_472 <= sw;
          th_myfunc_29 <= th_myfunc_29_6;
        end
        th_myfunc_29_6: begin
          _th_myfunc_29_i_473 <= 0;
          th_myfunc_29 <= th_myfunc_29_7;
        end
        th_myfunc_29_7: begin
          if(_th_myfunc_29_i_473 < _th_myfunc_29_time_472) begin
            th_myfunc_29 <= th_myfunc_29_8;
          end else begin
            th_myfunc_29 <= th_myfunc_29_12;
          end
        end
        th_myfunc_29_8: begin
          _th_myfunc_29___474 <= 0;
          th_myfunc_29 <= th_myfunc_29_9;
        end
        th_myfunc_29_9: begin
          if(_th_myfunc_29___474 < 1024) begin
            th_myfunc_29 <= th_myfunc_29_10;
          end else begin
            th_myfunc_29 <= th_myfunc_29_11;
          end
        end
        th_myfunc_29_10: begin
          _th_myfunc_29___474 <= _th_myfunc_29___474 + 1;
          th_myfunc_29 <= th_myfunc_29_9;
        end
        th_myfunc_29_11: begin
          _th_myfunc_29_i_473 <= _th_myfunc_29_i_473 + 1;
          th_myfunc_29 <= th_myfunc_29_7;
        end
        th_myfunc_29_12: begin
          th_myfunc_29 <= th_myfunc_29_13;
        end
        th_myfunc_29_13: begin
          $display("Thread %d count = %d", _th_myfunc_29_tid_471, count);
          th_myfunc_29 <= th_myfunc_29_14;
        end
        th_myfunc_29_14: begin
          th_myfunc_29 <= th_myfunc_29_15;
        end
        th_myfunc_29_15: begin
          $display("Thread %d Unlock", _th_myfunc_29_tid_471);
          th_myfunc_29 <= th_myfunc_29_16;
        end
        th_myfunc_29_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 29)) begin
            _th_myfunc_29_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 29)) begin
            th_myfunc_29 <= th_myfunc_29_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_30_1 = 1;
  localparam th_myfunc_30_2 = 2;
  localparam th_myfunc_30_3 = 3;
  localparam th_myfunc_30_4 = 4;
  localparam th_myfunc_30_5 = 5;
  localparam th_myfunc_30_6 = 6;
  localparam th_myfunc_30_7 = 7;
  localparam th_myfunc_30_8 = 8;
  localparam th_myfunc_30_9 = 9;
  localparam th_myfunc_30_10 = 10;
  localparam th_myfunc_30_11 = 11;
  localparam th_myfunc_30_12 = 12;
  localparam th_myfunc_30_13 = 13;
  localparam th_myfunc_30_14 = 14;
  localparam th_myfunc_30_15 = 15;
  localparam th_myfunc_30_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_30 <= th_myfunc_30_init;
      _th_myfunc_30_called <= 0;
      _th_myfunc_30_tid_475 <= 0;
      _th_myfunc_30_tid_476 <= 0;
      _th_myfunc_30_time_477 <= 0;
      _th_myfunc_30_i_478 <= 0;
      _th_myfunc_30___479 <= 0;
    end else begin
      case(th_myfunc_30)
        th_myfunc_30_init: begin
          if(_th_myfunc_start[30] && (th_blink == 10)) begin
            _th_myfunc_30_called <= 1;
          end 
          if(_th_myfunc_start[30] && (th_blink == 10)) begin
            _th_myfunc_30_tid_475 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[30]) begin
            th_myfunc_30 <= th_myfunc_30_1;
          end 
        end
        th_myfunc_30_1: begin
          _th_myfunc_30_tid_476 <= _th_myfunc_30_tid_475;
          th_myfunc_30 <= th_myfunc_30_2;
        end
        th_myfunc_30_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 30)) begin
            th_myfunc_30 <= th_myfunc_30_3;
          end 
        end
        th_myfunc_30_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 30))) begin
            th_myfunc_30 <= th_myfunc_30_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 30)) begin
            th_myfunc_30 <= th_myfunc_30_4;
          end 
        end
        th_myfunc_30_4: begin
          $display("Thread %d Lock", _th_myfunc_30_tid_476);
          th_myfunc_30 <= th_myfunc_30_5;
        end
        th_myfunc_30_5: begin
          _th_myfunc_30_time_477 <= sw;
          th_myfunc_30 <= th_myfunc_30_6;
        end
        th_myfunc_30_6: begin
          _th_myfunc_30_i_478 <= 0;
          th_myfunc_30 <= th_myfunc_30_7;
        end
        th_myfunc_30_7: begin
          if(_th_myfunc_30_i_478 < _th_myfunc_30_time_477) begin
            th_myfunc_30 <= th_myfunc_30_8;
          end else begin
            th_myfunc_30 <= th_myfunc_30_12;
          end
        end
        th_myfunc_30_8: begin
          _th_myfunc_30___479 <= 0;
          th_myfunc_30 <= th_myfunc_30_9;
        end
        th_myfunc_30_9: begin
          if(_th_myfunc_30___479 < 1024) begin
            th_myfunc_30 <= th_myfunc_30_10;
          end else begin
            th_myfunc_30 <= th_myfunc_30_11;
          end
        end
        th_myfunc_30_10: begin
          _th_myfunc_30___479 <= _th_myfunc_30___479 + 1;
          th_myfunc_30 <= th_myfunc_30_9;
        end
        th_myfunc_30_11: begin
          _th_myfunc_30_i_478 <= _th_myfunc_30_i_478 + 1;
          th_myfunc_30 <= th_myfunc_30_7;
        end
        th_myfunc_30_12: begin
          th_myfunc_30 <= th_myfunc_30_13;
        end
        th_myfunc_30_13: begin
          $display("Thread %d count = %d", _th_myfunc_30_tid_476, count);
          th_myfunc_30 <= th_myfunc_30_14;
        end
        th_myfunc_30_14: begin
          th_myfunc_30 <= th_myfunc_30_15;
        end
        th_myfunc_30_15: begin
          $display("Thread %d Unlock", _th_myfunc_30_tid_476);
          th_myfunc_30 <= th_myfunc_30_16;
        end
        th_myfunc_30_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 30)) begin
            _th_myfunc_30_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 30)) begin
            th_myfunc_30 <= th_myfunc_30_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_31_1 = 1;
  localparam th_myfunc_31_2 = 2;
  localparam th_myfunc_31_3 = 3;
  localparam th_myfunc_31_4 = 4;
  localparam th_myfunc_31_5 = 5;
  localparam th_myfunc_31_6 = 6;
  localparam th_myfunc_31_7 = 7;
  localparam th_myfunc_31_8 = 8;
  localparam th_myfunc_31_9 = 9;
  localparam th_myfunc_31_10 = 10;
  localparam th_myfunc_31_11 = 11;
  localparam th_myfunc_31_12 = 12;
  localparam th_myfunc_31_13 = 13;
  localparam th_myfunc_31_14 = 14;
  localparam th_myfunc_31_15 = 15;
  localparam th_myfunc_31_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_31 <= th_myfunc_31_init;
      _th_myfunc_31_called <= 0;
      _th_myfunc_31_tid_480 <= 0;
      _th_myfunc_31_tid_481 <= 0;
      _th_myfunc_31_time_482 <= 0;
      _th_myfunc_31_i_483 <= 0;
      _th_myfunc_31___484 <= 0;
    end else begin
      case(th_myfunc_31)
        th_myfunc_31_init: begin
          if(_th_myfunc_start[31] && (th_blink == 10)) begin
            _th_myfunc_31_called <= 1;
          end 
          if(_th_myfunc_start[31] && (th_blink == 10)) begin
            _th_myfunc_31_tid_480 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[31]) begin
            th_myfunc_31 <= th_myfunc_31_1;
          end 
        end
        th_myfunc_31_1: begin
          _th_myfunc_31_tid_481 <= _th_myfunc_31_tid_480;
          th_myfunc_31 <= th_myfunc_31_2;
        end
        th_myfunc_31_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 31)) begin
            th_myfunc_31 <= th_myfunc_31_3;
          end 
        end
        th_myfunc_31_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 31))) begin
            th_myfunc_31 <= th_myfunc_31_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 31)) begin
            th_myfunc_31 <= th_myfunc_31_4;
          end 
        end
        th_myfunc_31_4: begin
          $display("Thread %d Lock", _th_myfunc_31_tid_481);
          th_myfunc_31 <= th_myfunc_31_5;
        end
        th_myfunc_31_5: begin
          _th_myfunc_31_time_482 <= sw;
          th_myfunc_31 <= th_myfunc_31_6;
        end
        th_myfunc_31_6: begin
          _th_myfunc_31_i_483 <= 0;
          th_myfunc_31 <= th_myfunc_31_7;
        end
        th_myfunc_31_7: begin
          if(_th_myfunc_31_i_483 < _th_myfunc_31_time_482) begin
            th_myfunc_31 <= th_myfunc_31_8;
          end else begin
            th_myfunc_31 <= th_myfunc_31_12;
          end
        end
        th_myfunc_31_8: begin
          _th_myfunc_31___484 <= 0;
          th_myfunc_31 <= th_myfunc_31_9;
        end
        th_myfunc_31_9: begin
          if(_th_myfunc_31___484 < 1024) begin
            th_myfunc_31 <= th_myfunc_31_10;
          end else begin
            th_myfunc_31 <= th_myfunc_31_11;
          end
        end
        th_myfunc_31_10: begin
          _th_myfunc_31___484 <= _th_myfunc_31___484 + 1;
          th_myfunc_31 <= th_myfunc_31_9;
        end
        th_myfunc_31_11: begin
          _th_myfunc_31_i_483 <= _th_myfunc_31_i_483 + 1;
          th_myfunc_31 <= th_myfunc_31_7;
        end
        th_myfunc_31_12: begin
          th_myfunc_31 <= th_myfunc_31_13;
        end
        th_myfunc_31_13: begin
          $display("Thread %d count = %d", _th_myfunc_31_tid_481, count);
          th_myfunc_31 <= th_myfunc_31_14;
        end
        th_myfunc_31_14: begin
          th_myfunc_31 <= th_myfunc_31_15;
        end
        th_myfunc_31_15: begin
          $display("Thread %d Unlock", _th_myfunc_31_tid_481);
          th_myfunc_31 <= th_myfunc_31_16;
        end
        th_myfunc_31_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 31)) begin
            _th_myfunc_31_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 31)) begin
            th_myfunc_31 <= th_myfunc_31_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_32_1 = 1;
  localparam th_myfunc_32_2 = 2;
  localparam th_myfunc_32_3 = 3;
  localparam th_myfunc_32_4 = 4;
  localparam th_myfunc_32_5 = 5;
  localparam th_myfunc_32_6 = 6;
  localparam th_myfunc_32_7 = 7;
  localparam th_myfunc_32_8 = 8;
  localparam th_myfunc_32_9 = 9;
  localparam th_myfunc_32_10 = 10;
  localparam th_myfunc_32_11 = 11;
  localparam th_myfunc_32_12 = 12;
  localparam th_myfunc_32_13 = 13;
  localparam th_myfunc_32_14 = 14;
  localparam th_myfunc_32_15 = 15;
  localparam th_myfunc_32_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_32 <= th_myfunc_32_init;
      _th_myfunc_32_called <= 0;
      _th_myfunc_32_tid_485 <= 0;
      _th_myfunc_32_tid_486 <= 0;
      _th_myfunc_32_time_487 <= 0;
      _th_myfunc_32_i_488 <= 0;
      _th_myfunc_32___489 <= 0;
    end else begin
      case(th_myfunc_32)
        th_myfunc_32_init: begin
          if(_th_myfunc_start[32] && (th_blink == 10)) begin
            _th_myfunc_32_called <= 1;
          end 
          if(_th_myfunc_start[32] && (th_blink == 10)) begin
            _th_myfunc_32_tid_485 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[32]) begin
            th_myfunc_32 <= th_myfunc_32_1;
          end 
        end
        th_myfunc_32_1: begin
          _th_myfunc_32_tid_486 <= _th_myfunc_32_tid_485;
          th_myfunc_32 <= th_myfunc_32_2;
        end
        th_myfunc_32_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 32)) begin
            th_myfunc_32 <= th_myfunc_32_3;
          end 
        end
        th_myfunc_32_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 32))) begin
            th_myfunc_32 <= th_myfunc_32_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 32)) begin
            th_myfunc_32 <= th_myfunc_32_4;
          end 
        end
        th_myfunc_32_4: begin
          $display("Thread %d Lock", _th_myfunc_32_tid_486);
          th_myfunc_32 <= th_myfunc_32_5;
        end
        th_myfunc_32_5: begin
          _th_myfunc_32_time_487 <= sw;
          th_myfunc_32 <= th_myfunc_32_6;
        end
        th_myfunc_32_6: begin
          _th_myfunc_32_i_488 <= 0;
          th_myfunc_32 <= th_myfunc_32_7;
        end
        th_myfunc_32_7: begin
          if(_th_myfunc_32_i_488 < _th_myfunc_32_time_487) begin
            th_myfunc_32 <= th_myfunc_32_8;
          end else begin
            th_myfunc_32 <= th_myfunc_32_12;
          end
        end
        th_myfunc_32_8: begin
          _th_myfunc_32___489 <= 0;
          th_myfunc_32 <= th_myfunc_32_9;
        end
        th_myfunc_32_9: begin
          if(_th_myfunc_32___489 < 1024) begin
            th_myfunc_32 <= th_myfunc_32_10;
          end else begin
            th_myfunc_32 <= th_myfunc_32_11;
          end
        end
        th_myfunc_32_10: begin
          _th_myfunc_32___489 <= _th_myfunc_32___489 + 1;
          th_myfunc_32 <= th_myfunc_32_9;
        end
        th_myfunc_32_11: begin
          _th_myfunc_32_i_488 <= _th_myfunc_32_i_488 + 1;
          th_myfunc_32 <= th_myfunc_32_7;
        end
        th_myfunc_32_12: begin
          th_myfunc_32 <= th_myfunc_32_13;
        end
        th_myfunc_32_13: begin
          $display("Thread %d count = %d", _th_myfunc_32_tid_486, count);
          th_myfunc_32 <= th_myfunc_32_14;
        end
        th_myfunc_32_14: begin
          th_myfunc_32 <= th_myfunc_32_15;
        end
        th_myfunc_32_15: begin
          $display("Thread %d Unlock", _th_myfunc_32_tid_486);
          th_myfunc_32 <= th_myfunc_32_16;
        end
        th_myfunc_32_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 32)) begin
            _th_myfunc_32_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 32)) begin
            th_myfunc_32 <= th_myfunc_32_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_33_1 = 1;
  localparam th_myfunc_33_2 = 2;
  localparam th_myfunc_33_3 = 3;
  localparam th_myfunc_33_4 = 4;
  localparam th_myfunc_33_5 = 5;
  localparam th_myfunc_33_6 = 6;
  localparam th_myfunc_33_7 = 7;
  localparam th_myfunc_33_8 = 8;
  localparam th_myfunc_33_9 = 9;
  localparam th_myfunc_33_10 = 10;
  localparam th_myfunc_33_11 = 11;
  localparam th_myfunc_33_12 = 12;
  localparam th_myfunc_33_13 = 13;
  localparam th_myfunc_33_14 = 14;
  localparam th_myfunc_33_15 = 15;
  localparam th_myfunc_33_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_33 <= th_myfunc_33_init;
      _th_myfunc_33_called <= 0;
      _th_myfunc_33_tid_490 <= 0;
      _th_myfunc_33_tid_491 <= 0;
      _th_myfunc_33_time_492 <= 0;
      _th_myfunc_33_i_493 <= 0;
      _th_myfunc_33___494 <= 0;
    end else begin
      case(th_myfunc_33)
        th_myfunc_33_init: begin
          if(_th_myfunc_start[33] && (th_blink == 10)) begin
            _th_myfunc_33_called <= 1;
          end 
          if(_th_myfunc_start[33] && (th_blink == 10)) begin
            _th_myfunc_33_tid_490 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[33]) begin
            th_myfunc_33 <= th_myfunc_33_1;
          end 
        end
        th_myfunc_33_1: begin
          _th_myfunc_33_tid_491 <= _th_myfunc_33_tid_490;
          th_myfunc_33 <= th_myfunc_33_2;
        end
        th_myfunc_33_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 33)) begin
            th_myfunc_33 <= th_myfunc_33_3;
          end 
        end
        th_myfunc_33_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 33))) begin
            th_myfunc_33 <= th_myfunc_33_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 33)) begin
            th_myfunc_33 <= th_myfunc_33_4;
          end 
        end
        th_myfunc_33_4: begin
          $display("Thread %d Lock", _th_myfunc_33_tid_491);
          th_myfunc_33 <= th_myfunc_33_5;
        end
        th_myfunc_33_5: begin
          _th_myfunc_33_time_492 <= sw;
          th_myfunc_33 <= th_myfunc_33_6;
        end
        th_myfunc_33_6: begin
          _th_myfunc_33_i_493 <= 0;
          th_myfunc_33 <= th_myfunc_33_7;
        end
        th_myfunc_33_7: begin
          if(_th_myfunc_33_i_493 < _th_myfunc_33_time_492) begin
            th_myfunc_33 <= th_myfunc_33_8;
          end else begin
            th_myfunc_33 <= th_myfunc_33_12;
          end
        end
        th_myfunc_33_8: begin
          _th_myfunc_33___494 <= 0;
          th_myfunc_33 <= th_myfunc_33_9;
        end
        th_myfunc_33_9: begin
          if(_th_myfunc_33___494 < 1024) begin
            th_myfunc_33 <= th_myfunc_33_10;
          end else begin
            th_myfunc_33 <= th_myfunc_33_11;
          end
        end
        th_myfunc_33_10: begin
          _th_myfunc_33___494 <= _th_myfunc_33___494 + 1;
          th_myfunc_33 <= th_myfunc_33_9;
        end
        th_myfunc_33_11: begin
          _th_myfunc_33_i_493 <= _th_myfunc_33_i_493 + 1;
          th_myfunc_33 <= th_myfunc_33_7;
        end
        th_myfunc_33_12: begin
          th_myfunc_33 <= th_myfunc_33_13;
        end
        th_myfunc_33_13: begin
          $display("Thread %d count = %d", _th_myfunc_33_tid_491, count);
          th_myfunc_33 <= th_myfunc_33_14;
        end
        th_myfunc_33_14: begin
          th_myfunc_33 <= th_myfunc_33_15;
        end
        th_myfunc_33_15: begin
          $display("Thread %d Unlock", _th_myfunc_33_tid_491);
          th_myfunc_33 <= th_myfunc_33_16;
        end
        th_myfunc_33_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 33)) begin
            _th_myfunc_33_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 33)) begin
            th_myfunc_33 <= th_myfunc_33_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_34_1 = 1;
  localparam th_myfunc_34_2 = 2;
  localparam th_myfunc_34_3 = 3;
  localparam th_myfunc_34_4 = 4;
  localparam th_myfunc_34_5 = 5;
  localparam th_myfunc_34_6 = 6;
  localparam th_myfunc_34_7 = 7;
  localparam th_myfunc_34_8 = 8;
  localparam th_myfunc_34_9 = 9;
  localparam th_myfunc_34_10 = 10;
  localparam th_myfunc_34_11 = 11;
  localparam th_myfunc_34_12 = 12;
  localparam th_myfunc_34_13 = 13;
  localparam th_myfunc_34_14 = 14;
  localparam th_myfunc_34_15 = 15;
  localparam th_myfunc_34_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_34 <= th_myfunc_34_init;
      _th_myfunc_34_called <= 0;
      _th_myfunc_34_tid_495 <= 0;
      _th_myfunc_34_tid_496 <= 0;
      _th_myfunc_34_time_497 <= 0;
      _th_myfunc_34_i_498 <= 0;
      _th_myfunc_34___499 <= 0;
    end else begin
      case(th_myfunc_34)
        th_myfunc_34_init: begin
          if(_th_myfunc_start[34] && (th_blink == 10)) begin
            _th_myfunc_34_called <= 1;
          end 
          if(_th_myfunc_start[34] && (th_blink == 10)) begin
            _th_myfunc_34_tid_495 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[34]) begin
            th_myfunc_34 <= th_myfunc_34_1;
          end 
        end
        th_myfunc_34_1: begin
          _th_myfunc_34_tid_496 <= _th_myfunc_34_tid_495;
          th_myfunc_34 <= th_myfunc_34_2;
        end
        th_myfunc_34_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 34)) begin
            th_myfunc_34 <= th_myfunc_34_3;
          end 
        end
        th_myfunc_34_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 34))) begin
            th_myfunc_34 <= th_myfunc_34_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 34)) begin
            th_myfunc_34 <= th_myfunc_34_4;
          end 
        end
        th_myfunc_34_4: begin
          $display("Thread %d Lock", _th_myfunc_34_tid_496);
          th_myfunc_34 <= th_myfunc_34_5;
        end
        th_myfunc_34_5: begin
          _th_myfunc_34_time_497 <= sw;
          th_myfunc_34 <= th_myfunc_34_6;
        end
        th_myfunc_34_6: begin
          _th_myfunc_34_i_498 <= 0;
          th_myfunc_34 <= th_myfunc_34_7;
        end
        th_myfunc_34_7: begin
          if(_th_myfunc_34_i_498 < _th_myfunc_34_time_497) begin
            th_myfunc_34 <= th_myfunc_34_8;
          end else begin
            th_myfunc_34 <= th_myfunc_34_12;
          end
        end
        th_myfunc_34_8: begin
          _th_myfunc_34___499 <= 0;
          th_myfunc_34 <= th_myfunc_34_9;
        end
        th_myfunc_34_9: begin
          if(_th_myfunc_34___499 < 1024) begin
            th_myfunc_34 <= th_myfunc_34_10;
          end else begin
            th_myfunc_34 <= th_myfunc_34_11;
          end
        end
        th_myfunc_34_10: begin
          _th_myfunc_34___499 <= _th_myfunc_34___499 + 1;
          th_myfunc_34 <= th_myfunc_34_9;
        end
        th_myfunc_34_11: begin
          _th_myfunc_34_i_498 <= _th_myfunc_34_i_498 + 1;
          th_myfunc_34 <= th_myfunc_34_7;
        end
        th_myfunc_34_12: begin
          th_myfunc_34 <= th_myfunc_34_13;
        end
        th_myfunc_34_13: begin
          $display("Thread %d count = %d", _th_myfunc_34_tid_496, count);
          th_myfunc_34 <= th_myfunc_34_14;
        end
        th_myfunc_34_14: begin
          th_myfunc_34 <= th_myfunc_34_15;
        end
        th_myfunc_34_15: begin
          $display("Thread %d Unlock", _th_myfunc_34_tid_496);
          th_myfunc_34 <= th_myfunc_34_16;
        end
        th_myfunc_34_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 34)) begin
            _th_myfunc_34_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 34)) begin
            th_myfunc_34 <= th_myfunc_34_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_35_1 = 1;
  localparam th_myfunc_35_2 = 2;
  localparam th_myfunc_35_3 = 3;
  localparam th_myfunc_35_4 = 4;
  localparam th_myfunc_35_5 = 5;
  localparam th_myfunc_35_6 = 6;
  localparam th_myfunc_35_7 = 7;
  localparam th_myfunc_35_8 = 8;
  localparam th_myfunc_35_9 = 9;
  localparam th_myfunc_35_10 = 10;
  localparam th_myfunc_35_11 = 11;
  localparam th_myfunc_35_12 = 12;
  localparam th_myfunc_35_13 = 13;
  localparam th_myfunc_35_14 = 14;
  localparam th_myfunc_35_15 = 15;
  localparam th_myfunc_35_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_35 <= th_myfunc_35_init;
      _th_myfunc_35_called <= 0;
      _th_myfunc_35_tid_500 <= 0;
      _th_myfunc_35_tid_501 <= 0;
      _th_myfunc_35_time_502 <= 0;
      _th_myfunc_35_i_503 <= 0;
      _th_myfunc_35___504 <= 0;
    end else begin
      case(th_myfunc_35)
        th_myfunc_35_init: begin
          if(_th_myfunc_start[35] && (th_blink == 10)) begin
            _th_myfunc_35_called <= 1;
          end 
          if(_th_myfunc_start[35] && (th_blink == 10)) begin
            _th_myfunc_35_tid_500 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[35]) begin
            th_myfunc_35 <= th_myfunc_35_1;
          end 
        end
        th_myfunc_35_1: begin
          _th_myfunc_35_tid_501 <= _th_myfunc_35_tid_500;
          th_myfunc_35 <= th_myfunc_35_2;
        end
        th_myfunc_35_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 35)) begin
            th_myfunc_35 <= th_myfunc_35_3;
          end 
        end
        th_myfunc_35_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 35))) begin
            th_myfunc_35 <= th_myfunc_35_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 35)) begin
            th_myfunc_35 <= th_myfunc_35_4;
          end 
        end
        th_myfunc_35_4: begin
          $display("Thread %d Lock", _th_myfunc_35_tid_501);
          th_myfunc_35 <= th_myfunc_35_5;
        end
        th_myfunc_35_5: begin
          _th_myfunc_35_time_502 <= sw;
          th_myfunc_35 <= th_myfunc_35_6;
        end
        th_myfunc_35_6: begin
          _th_myfunc_35_i_503 <= 0;
          th_myfunc_35 <= th_myfunc_35_7;
        end
        th_myfunc_35_7: begin
          if(_th_myfunc_35_i_503 < _th_myfunc_35_time_502) begin
            th_myfunc_35 <= th_myfunc_35_8;
          end else begin
            th_myfunc_35 <= th_myfunc_35_12;
          end
        end
        th_myfunc_35_8: begin
          _th_myfunc_35___504 <= 0;
          th_myfunc_35 <= th_myfunc_35_9;
        end
        th_myfunc_35_9: begin
          if(_th_myfunc_35___504 < 1024) begin
            th_myfunc_35 <= th_myfunc_35_10;
          end else begin
            th_myfunc_35 <= th_myfunc_35_11;
          end
        end
        th_myfunc_35_10: begin
          _th_myfunc_35___504 <= _th_myfunc_35___504 + 1;
          th_myfunc_35 <= th_myfunc_35_9;
        end
        th_myfunc_35_11: begin
          _th_myfunc_35_i_503 <= _th_myfunc_35_i_503 + 1;
          th_myfunc_35 <= th_myfunc_35_7;
        end
        th_myfunc_35_12: begin
          th_myfunc_35 <= th_myfunc_35_13;
        end
        th_myfunc_35_13: begin
          $display("Thread %d count = %d", _th_myfunc_35_tid_501, count);
          th_myfunc_35 <= th_myfunc_35_14;
        end
        th_myfunc_35_14: begin
          th_myfunc_35 <= th_myfunc_35_15;
        end
        th_myfunc_35_15: begin
          $display("Thread %d Unlock", _th_myfunc_35_tid_501);
          th_myfunc_35 <= th_myfunc_35_16;
        end
        th_myfunc_35_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 35)) begin
            _th_myfunc_35_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 35)) begin
            th_myfunc_35 <= th_myfunc_35_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_36_1 = 1;
  localparam th_myfunc_36_2 = 2;
  localparam th_myfunc_36_3 = 3;
  localparam th_myfunc_36_4 = 4;
  localparam th_myfunc_36_5 = 5;
  localparam th_myfunc_36_6 = 6;
  localparam th_myfunc_36_7 = 7;
  localparam th_myfunc_36_8 = 8;
  localparam th_myfunc_36_9 = 9;
  localparam th_myfunc_36_10 = 10;
  localparam th_myfunc_36_11 = 11;
  localparam th_myfunc_36_12 = 12;
  localparam th_myfunc_36_13 = 13;
  localparam th_myfunc_36_14 = 14;
  localparam th_myfunc_36_15 = 15;
  localparam th_myfunc_36_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_36 <= th_myfunc_36_init;
      _th_myfunc_36_called <= 0;
      _th_myfunc_36_tid_505 <= 0;
      _th_myfunc_36_tid_506 <= 0;
      _th_myfunc_36_time_507 <= 0;
      _th_myfunc_36_i_508 <= 0;
      _th_myfunc_36___509 <= 0;
    end else begin
      case(th_myfunc_36)
        th_myfunc_36_init: begin
          if(_th_myfunc_start[36] && (th_blink == 10)) begin
            _th_myfunc_36_called <= 1;
          end 
          if(_th_myfunc_start[36] && (th_blink == 10)) begin
            _th_myfunc_36_tid_505 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[36]) begin
            th_myfunc_36 <= th_myfunc_36_1;
          end 
        end
        th_myfunc_36_1: begin
          _th_myfunc_36_tid_506 <= _th_myfunc_36_tid_505;
          th_myfunc_36 <= th_myfunc_36_2;
        end
        th_myfunc_36_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 36)) begin
            th_myfunc_36 <= th_myfunc_36_3;
          end 
        end
        th_myfunc_36_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 36))) begin
            th_myfunc_36 <= th_myfunc_36_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 36)) begin
            th_myfunc_36 <= th_myfunc_36_4;
          end 
        end
        th_myfunc_36_4: begin
          $display("Thread %d Lock", _th_myfunc_36_tid_506);
          th_myfunc_36 <= th_myfunc_36_5;
        end
        th_myfunc_36_5: begin
          _th_myfunc_36_time_507 <= sw;
          th_myfunc_36 <= th_myfunc_36_6;
        end
        th_myfunc_36_6: begin
          _th_myfunc_36_i_508 <= 0;
          th_myfunc_36 <= th_myfunc_36_7;
        end
        th_myfunc_36_7: begin
          if(_th_myfunc_36_i_508 < _th_myfunc_36_time_507) begin
            th_myfunc_36 <= th_myfunc_36_8;
          end else begin
            th_myfunc_36 <= th_myfunc_36_12;
          end
        end
        th_myfunc_36_8: begin
          _th_myfunc_36___509 <= 0;
          th_myfunc_36 <= th_myfunc_36_9;
        end
        th_myfunc_36_9: begin
          if(_th_myfunc_36___509 < 1024) begin
            th_myfunc_36 <= th_myfunc_36_10;
          end else begin
            th_myfunc_36 <= th_myfunc_36_11;
          end
        end
        th_myfunc_36_10: begin
          _th_myfunc_36___509 <= _th_myfunc_36___509 + 1;
          th_myfunc_36 <= th_myfunc_36_9;
        end
        th_myfunc_36_11: begin
          _th_myfunc_36_i_508 <= _th_myfunc_36_i_508 + 1;
          th_myfunc_36 <= th_myfunc_36_7;
        end
        th_myfunc_36_12: begin
          th_myfunc_36 <= th_myfunc_36_13;
        end
        th_myfunc_36_13: begin
          $display("Thread %d count = %d", _th_myfunc_36_tid_506, count);
          th_myfunc_36 <= th_myfunc_36_14;
        end
        th_myfunc_36_14: begin
          th_myfunc_36 <= th_myfunc_36_15;
        end
        th_myfunc_36_15: begin
          $display("Thread %d Unlock", _th_myfunc_36_tid_506);
          th_myfunc_36 <= th_myfunc_36_16;
        end
        th_myfunc_36_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 36)) begin
            _th_myfunc_36_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 36)) begin
            th_myfunc_36 <= th_myfunc_36_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_37_1 = 1;
  localparam th_myfunc_37_2 = 2;
  localparam th_myfunc_37_3 = 3;
  localparam th_myfunc_37_4 = 4;
  localparam th_myfunc_37_5 = 5;
  localparam th_myfunc_37_6 = 6;
  localparam th_myfunc_37_7 = 7;
  localparam th_myfunc_37_8 = 8;
  localparam th_myfunc_37_9 = 9;
  localparam th_myfunc_37_10 = 10;
  localparam th_myfunc_37_11 = 11;
  localparam th_myfunc_37_12 = 12;
  localparam th_myfunc_37_13 = 13;
  localparam th_myfunc_37_14 = 14;
  localparam th_myfunc_37_15 = 15;
  localparam th_myfunc_37_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_37 <= th_myfunc_37_init;
      _th_myfunc_37_called <= 0;
      _th_myfunc_37_tid_510 <= 0;
      _th_myfunc_37_tid_511 <= 0;
      _th_myfunc_37_time_512 <= 0;
      _th_myfunc_37_i_513 <= 0;
      _th_myfunc_37___514 <= 0;
    end else begin
      case(th_myfunc_37)
        th_myfunc_37_init: begin
          if(_th_myfunc_start[37] && (th_blink == 10)) begin
            _th_myfunc_37_called <= 1;
          end 
          if(_th_myfunc_start[37] && (th_blink == 10)) begin
            _th_myfunc_37_tid_510 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[37]) begin
            th_myfunc_37 <= th_myfunc_37_1;
          end 
        end
        th_myfunc_37_1: begin
          _th_myfunc_37_tid_511 <= _th_myfunc_37_tid_510;
          th_myfunc_37 <= th_myfunc_37_2;
        end
        th_myfunc_37_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 37)) begin
            th_myfunc_37 <= th_myfunc_37_3;
          end 
        end
        th_myfunc_37_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 37))) begin
            th_myfunc_37 <= th_myfunc_37_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 37)) begin
            th_myfunc_37 <= th_myfunc_37_4;
          end 
        end
        th_myfunc_37_4: begin
          $display("Thread %d Lock", _th_myfunc_37_tid_511);
          th_myfunc_37 <= th_myfunc_37_5;
        end
        th_myfunc_37_5: begin
          _th_myfunc_37_time_512 <= sw;
          th_myfunc_37 <= th_myfunc_37_6;
        end
        th_myfunc_37_6: begin
          _th_myfunc_37_i_513 <= 0;
          th_myfunc_37 <= th_myfunc_37_7;
        end
        th_myfunc_37_7: begin
          if(_th_myfunc_37_i_513 < _th_myfunc_37_time_512) begin
            th_myfunc_37 <= th_myfunc_37_8;
          end else begin
            th_myfunc_37 <= th_myfunc_37_12;
          end
        end
        th_myfunc_37_8: begin
          _th_myfunc_37___514 <= 0;
          th_myfunc_37 <= th_myfunc_37_9;
        end
        th_myfunc_37_9: begin
          if(_th_myfunc_37___514 < 1024) begin
            th_myfunc_37 <= th_myfunc_37_10;
          end else begin
            th_myfunc_37 <= th_myfunc_37_11;
          end
        end
        th_myfunc_37_10: begin
          _th_myfunc_37___514 <= _th_myfunc_37___514 + 1;
          th_myfunc_37 <= th_myfunc_37_9;
        end
        th_myfunc_37_11: begin
          _th_myfunc_37_i_513 <= _th_myfunc_37_i_513 + 1;
          th_myfunc_37 <= th_myfunc_37_7;
        end
        th_myfunc_37_12: begin
          th_myfunc_37 <= th_myfunc_37_13;
        end
        th_myfunc_37_13: begin
          $display("Thread %d count = %d", _th_myfunc_37_tid_511, count);
          th_myfunc_37 <= th_myfunc_37_14;
        end
        th_myfunc_37_14: begin
          th_myfunc_37 <= th_myfunc_37_15;
        end
        th_myfunc_37_15: begin
          $display("Thread %d Unlock", _th_myfunc_37_tid_511);
          th_myfunc_37 <= th_myfunc_37_16;
        end
        th_myfunc_37_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 37)) begin
            _th_myfunc_37_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 37)) begin
            th_myfunc_37 <= th_myfunc_37_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_38_1 = 1;
  localparam th_myfunc_38_2 = 2;
  localparam th_myfunc_38_3 = 3;
  localparam th_myfunc_38_4 = 4;
  localparam th_myfunc_38_5 = 5;
  localparam th_myfunc_38_6 = 6;
  localparam th_myfunc_38_7 = 7;
  localparam th_myfunc_38_8 = 8;
  localparam th_myfunc_38_9 = 9;
  localparam th_myfunc_38_10 = 10;
  localparam th_myfunc_38_11 = 11;
  localparam th_myfunc_38_12 = 12;
  localparam th_myfunc_38_13 = 13;
  localparam th_myfunc_38_14 = 14;
  localparam th_myfunc_38_15 = 15;
  localparam th_myfunc_38_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_38 <= th_myfunc_38_init;
      _th_myfunc_38_called <= 0;
      _th_myfunc_38_tid_515 <= 0;
      _th_myfunc_38_tid_516 <= 0;
      _th_myfunc_38_time_517 <= 0;
      _th_myfunc_38_i_518 <= 0;
      _th_myfunc_38___519 <= 0;
    end else begin
      case(th_myfunc_38)
        th_myfunc_38_init: begin
          if(_th_myfunc_start[38] && (th_blink == 10)) begin
            _th_myfunc_38_called <= 1;
          end 
          if(_th_myfunc_start[38] && (th_blink == 10)) begin
            _th_myfunc_38_tid_515 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[38]) begin
            th_myfunc_38 <= th_myfunc_38_1;
          end 
        end
        th_myfunc_38_1: begin
          _th_myfunc_38_tid_516 <= _th_myfunc_38_tid_515;
          th_myfunc_38 <= th_myfunc_38_2;
        end
        th_myfunc_38_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 38)) begin
            th_myfunc_38 <= th_myfunc_38_3;
          end 
        end
        th_myfunc_38_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 38))) begin
            th_myfunc_38 <= th_myfunc_38_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 38)) begin
            th_myfunc_38 <= th_myfunc_38_4;
          end 
        end
        th_myfunc_38_4: begin
          $display("Thread %d Lock", _th_myfunc_38_tid_516);
          th_myfunc_38 <= th_myfunc_38_5;
        end
        th_myfunc_38_5: begin
          _th_myfunc_38_time_517 <= sw;
          th_myfunc_38 <= th_myfunc_38_6;
        end
        th_myfunc_38_6: begin
          _th_myfunc_38_i_518 <= 0;
          th_myfunc_38 <= th_myfunc_38_7;
        end
        th_myfunc_38_7: begin
          if(_th_myfunc_38_i_518 < _th_myfunc_38_time_517) begin
            th_myfunc_38 <= th_myfunc_38_8;
          end else begin
            th_myfunc_38 <= th_myfunc_38_12;
          end
        end
        th_myfunc_38_8: begin
          _th_myfunc_38___519 <= 0;
          th_myfunc_38 <= th_myfunc_38_9;
        end
        th_myfunc_38_9: begin
          if(_th_myfunc_38___519 < 1024) begin
            th_myfunc_38 <= th_myfunc_38_10;
          end else begin
            th_myfunc_38 <= th_myfunc_38_11;
          end
        end
        th_myfunc_38_10: begin
          _th_myfunc_38___519 <= _th_myfunc_38___519 + 1;
          th_myfunc_38 <= th_myfunc_38_9;
        end
        th_myfunc_38_11: begin
          _th_myfunc_38_i_518 <= _th_myfunc_38_i_518 + 1;
          th_myfunc_38 <= th_myfunc_38_7;
        end
        th_myfunc_38_12: begin
          th_myfunc_38 <= th_myfunc_38_13;
        end
        th_myfunc_38_13: begin
          $display("Thread %d count = %d", _th_myfunc_38_tid_516, count);
          th_myfunc_38 <= th_myfunc_38_14;
        end
        th_myfunc_38_14: begin
          th_myfunc_38 <= th_myfunc_38_15;
        end
        th_myfunc_38_15: begin
          $display("Thread %d Unlock", _th_myfunc_38_tid_516);
          th_myfunc_38 <= th_myfunc_38_16;
        end
        th_myfunc_38_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 38)) begin
            _th_myfunc_38_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 38)) begin
            th_myfunc_38 <= th_myfunc_38_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_39_1 = 1;
  localparam th_myfunc_39_2 = 2;
  localparam th_myfunc_39_3 = 3;
  localparam th_myfunc_39_4 = 4;
  localparam th_myfunc_39_5 = 5;
  localparam th_myfunc_39_6 = 6;
  localparam th_myfunc_39_7 = 7;
  localparam th_myfunc_39_8 = 8;
  localparam th_myfunc_39_9 = 9;
  localparam th_myfunc_39_10 = 10;
  localparam th_myfunc_39_11 = 11;
  localparam th_myfunc_39_12 = 12;
  localparam th_myfunc_39_13 = 13;
  localparam th_myfunc_39_14 = 14;
  localparam th_myfunc_39_15 = 15;
  localparam th_myfunc_39_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_39 <= th_myfunc_39_init;
      _th_myfunc_39_called <= 0;
      _th_myfunc_39_tid_520 <= 0;
      _th_myfunc_39_tid_521 <= 0;
      _th_myfunc_39_time_522 <= 0;
      _th_myfunc_39_i_523 <= 0;
      _th_myfunc_39___524 <= 0;
    end else begin
      case(th_myfunc_39)
        th_myfunc_39_init: begin
          if(_th_myfunc_start[39] && (th_blink == 10)) begin
            _th_myfunc_39_called <= 1;
          end 
          if(_th_myfunc_start[39] && (th_blink == 10)) begin
            _th_myfunc_39_tid_520 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[39]) begin
            th_myfunc_39 <= th_myfunc_39_1;
          end 
        end
        th_myfunc_39_1: begin
          _th_myfunc_39_tid_521 <= _th_myfunc_39_tid_520;
          th_myfunc_39 <= th_myfunc_39_2;
        end
        th_myfunc_39_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 39)) begin
            th_myfunc_39 <= th_myfunc_39_3;
          end 
        end
        th_myfunc_39_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 39))) begin
            th_myfunc_39 <= th_myfunc_39_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 39)) begin
            th_myfunc_39 <= th_myfunc_39_4;
          end 
        end
        th_myfunc_39_4: begin
          $display("Thread %d Lock", _th_myfunc_39_tid_521);
          th_myfunc_39 <= th_myfunc_39_5;
        end
        th_myfunc_39_5: begin
          _th_myfunc_39_time_522 <= sw;
          th_myfunc_39 <= th_myfunc_39_6;
        end
        th_myfunc_39_6: begin
          _th_myfunc_39_i_523 <= 0;
          th_myfunc_39 <= th_myfunc_39_7;
        end
        th_myfunc_39_7: begin
          if(_th_myfunc_39_i_523 < _th_myfunc_39_time_522) begin
            th_myfunc_39 <= th_myfunc_39_8;
          end else begin
            th_myfunc_39 <= th_myfunc_39_12;
          end
        end
        th_myfunc_39_8: begin
          _th_myfunc_39___524 <= 0;
          th_myfunc_39 <= th_myfunc_39_9;
        end
        th_myfunc_39_9: begin
          if(_th_myfunc_39___524 < 1024) begin
            th_myfunc_39 <= th_myfunc_39_10;
          end else begin
            th_myfunc_39 <= th_myfunc_39_11;
          end
        end
        th_myfunc_39_10: begin
          _th_myfunc_39___524 <= _th_myfunc_39___524 + 1;
          th_myfunc_39 <= th_myfunc_39_9;
        end
        th_myfunc_39_11: begin
          _th_myfunc_39_i_523 <= _th_myfunc_39_i_523 + 1;
          th_myfunc_39 <= th_myfunc_39_7;
        end
        th_myfunc_39_12: begin
          th_myfunc_39 <= th_myfunc_39_13;
        end
        th_myfunc_39_13: begin
          $display("Thread %d count = %d", _th_myfunc_39_tid_521, count);
          th_myfunc_39 <= th_myfunc_39_14;
        end
        th_myfunc_39_14: begin
          th_myfunc_39 <= th_myfunc_39_15;
        end
        th_myfunc_39_15: begin
          $display("Thread %d Unlock", _th_myfunc_39_tid_521);
          th_myfunc_39 <= th_myfunc_39_16;
        end
        th_myfunc_39_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 39)) begin
            _th_myfunc_39_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 39)) begin
            th_myfunc_39 <= th_myfunc_39_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_40_1 = 1;
  localparam th_myfunc_40_2 = 2;
  localparam th_myfunc_40_3 = 3;
  localparam th_myfunc_40_4 = 4;
  localparam th_myfunc_40_5 = 5;
  localparam th_myfunc_40_6 = 6;
  localparam th_myfunc_40_7 = 7;
  localparam th_myfunc_40_8 = 8;
  localparam th_myfunc_40_9 = 9;
  localparam th_myfunc_40_10 = 10;
  localparam th_myfunc_40_11 = 11;
  localparam th_myfunc_40_12 = 12;
  localparam th_myfunc_40_13 = 13;
  localparam th_myfunc_40_14 = 14;
  localparam th_myfunc_40_15 = 15;
  localparam th_myfunc_40_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_40 <= th_myfunc_40_init;
      _th_myfunc_40_called <= 0;
      _th_myfunc_40_tid_525 <= 0;
      _th_myfunc_40_tid_526 <= 0;
      _th_myfunc_40_time_527 <= 0;
      _th_myfunc_40_i_528 <= 0;
      _th_myfunc_40___529 <= 0;
    end else begin
      case(th_myfunc_40)
        th_myfunc_40_init: begin
          if(_th_myfunc_start[40] && (th_blink == 10)) begin
            _th_myfunc_40_called <= 1;
          end 
          if(_th_myfunc_start[40] && (th_blink == 10)) begin
            _th_myfunc_40_tid_525 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[40]) begin
            th_myfunc_40 <= th_myfunc_40_1;
          end 
        end
        th_myfunc_40_1: begin
          _th_myfunc_40_tid_526 <= _th_myfunc_40_tid_525;
          th_myfunc_40 <= th_myfunc_40_2;
        end
        th_myfunc_40_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 40)) begin
            th_myfunc_40 <= th_myfunc_40_3;
          end 
        end
        th_myfunc_40_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 40))) begin
            th_myfunc_40 <= th_myfunc_40_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 40)) begin
            th_myfunc_40 <= th_myfunc_40_4;
          end 
        end
        th_myfunc_40_4: begin
          $display("Thread %d Lock", _th_myfunc_40_tid_526);
          th_myfunc_40 <= th_myfunc_40_5;
        end
        th_myfunc_40_5: begin
          _th_myfunc_40_time_527 <= sw;
          th_myfunc_40 <= th_myfunc_40_6;
        end
        th_myfunc_40_6: begin
          _th_myfunc_40_i_528 <= 0;
          th_myfunc_40 <= th_myfunc_40_7;
        end
        th_myfunc_40_7: begin
          if(_th_myfunc_40_i_528 < _th_myfunc_40_time_527) begin
            th_myfunc_40 <= th_myfunc_40_8;
          end else begin
            th_myfunc_40 <= th_myfunc_40_12;
          end
        end
        th_myfunc_40_8: begin
          _th_myfunc_40___529 <= 0;
          th_myfunc_40 <= th_myfunc_40_9;
        end
        th_myfunc_40_9: begin
          if(_th_myfunc_40___529 < 1024) begin
            th_myfunc_40 <= th_myfunc_40_10;
          end else begin
            th_myfunc_40 <= th_myfunc_40_11;
          end
        end
        th_myfunc_40_10: begin
          _th_myfunc_40___529 <= _th_myfunc_40___529 + 1;
          th_myfunc_40 <= th_myfunc_40_9;
        end
        th_myfunc_40_11: begin
          _th_myfunc_40_i_528 <= _th_myfunc_40_i_528 + 1;
          th_myfunc_40 <= th_myfunc_40_7;
        end
        th_myfunc_40_12: begin
          th_myfunc_40 <= th_myfunc_40_13;
        end
        th_myfunc_40_13: begin
          $display("Thread %d count = %d", _th_myfunc_40_tid_526, count);
          th_myfunc_40 <= th_myfunc_40_14;
        end
        th_myfunc_40_14: begin
          th_myfunc_40 <= th_myfunc_40_15;
        end
        th_myfunc_40_15: begin
          $display("Thread %d Unlock", _th_myfunc_40_tid_526);
          th_myfunc_40 <= th_myfunc_40_16;
        end
        th_myfunc_40_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 40)) begin
            _th_myfunc_40_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 40)) begin
            th_myfunc_40 <= th_myfunc_40_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_41_1 = 1;
  localparam th_myfunc_41_2 = 2;
  localparam th_myfunc_41_3 = 3;
  localparam th_myfunc_41_4 = 4;
  localparam th_myfunc_41_5 = 5;
  localparam th_myfunc_41_6 = 6;
  localparam th_myfunc_41_7 = 7;
  localparam th_myfunc_41_8 = 8;
  localparam th_myfunc_41_9 = 9;
  localparam th_myfunc_41_10 = 10;
  localparam th_myfunc_41_11 = 11;
  localparam th_myfunc_41_12 = 12;
  localparam th_myfunc_41_13 = 13;
  localparam th_myfunc_41_14 = 14;
  localparam th_myfunc_41_15 = 15;
  localparam th_myfunc_41_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_41 <= th_myfunc_41_init;
      _th_myfunc_41_called <= 0;
      _th_myfunc_41_tid_530 <= 0;
      _th_myfunc_41_tid_531 <= 0;
      _th_myfunc_41_time_532 <= 0;
      _th_myfunc_41_i_533 <= 0;
      _th_myfunc_41___534 <= 0;
    end else begin
      case(th_myfunc_41)
        th_myfunc_41_init: begin
          if(_th_myfunc_start[41] && (th_blink == 10)) begin
            _th_myfunc_41_called <= 1;
          end 
          if(_th_myfunc_start[41] && (th_blink == 10)) begin
            _th_myfunc_41_tid_530 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[41]) begin
            th_myfunc_41 <= th_myfunc_41_1;
          end 
        end
        th_myfunc_41_1: begin
          _th_myfunc_41_tid_531 <= _th_myfunc_41_tid_530;
          th_myfunc_41 <= th_myfunc_41_2;
        end
        th_myfunc_41_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 41)) begin
            th_myfunc_41 <= th_myfunc_41_3;
          end 
        end
        th_myfunc_41_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 41))) begin
            th_myfunc_41 <= th_myfunc_41_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 41)) begin
            th_myfunc_41 <= th_myfunc_41_4;
          end 
        end
        th_myfunc_41_4: begin
          $display("Thread %d Lock", _th_myfunc_41_tid_531);
          th_myfunc_41 <= th_myfunc_41_5;
        end
        th_myfunc_41_5: begin
          _th_myfunc_41_time_532 <= sw;
          th_myfunc_41 <= th_myfunc_41_6;
        end
        th_myfunc_41_6: begin
          _th_myfunc_41_i_533 <= 0;
          th_myfunc_41 <= th_myfunc_41_7;
        end
        th_myfunc_41_7: begin
          if(_th_myfunc_41_i_533 < _th_myfunc_41_time_532) begin
            th_myfunc_41 <= th_myfunc_41_8;
          end else begin
            th_myfunc_41 <= th_myfunc_41_12;
          end
        end
        th_myfunc_41_8: begin
          _th_myfunc_41___534 <= 0;
          th_myfunc_41 <= th_myfunc_41_9;
        end
        th_myfunc_41_9: begin
          if(_th_myfunc_41___534 < 1024) begin
            th_myfunc_41 <= th_myfunc_41_10;
          end else begin
            th_myfunc_41 <= th_myfunc_41_11;
          end
        end
        th_myfunc_41_10: begin
          _th_myfunc_41___534 <= _th_myfunc_41___534 + 1;
          th_myfunc_41 <= th_myfunc_41_9;
        end
        th_myfunc_41_11: begin
          _th_myfunc_41_i_533 <= _th_myfunc_41_i_533 + 1;
          th_myfunc_41 <= th_myfunc_41_7;
        end
        th_myfunc_41_12: begin
          th_myfunc_41 <= th_myfunc_41_13;
        end
        th_myfunc_41_13: begin
          $display("Thread %d count = %d", _th_myfunc_41_tid_531, count);
          th_myfunc_41 <= th_myfunc_41_14;
        end
        th_myfunc_41_14: begin
          th_myfunc_41 <= th_myfunc_41_15;
        end
        th_myfunc_41_15: begin
          $display("Thread %d Unlock", _th_myfunc_41_tid_531);
          th_myfunc_41 <= th_myfunc_41_16;
        end
        th_myfunc_41_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 41)) begin
            _th_myfunc_41_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 41)) begin
            th_myfunc_41 <= th_myfunc_41_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_42_1 = 1;
  localparam th_myfunc_42_2 = 2;
  localparam th_myfunc_42_3 = 3;
  localparam th_myfunc_42_4 = 4;
  localparam th_myfunc_42_5 = 5;
  localparam th_myfunc_42_6 = 6;
  localparam th_myfunc_42_7 = 7;
  localparam th_myfunc_42_8 = 8;
  localparam th_myfunc_42_9 = 9;
  localparam th_myfunc_42_10 = 10;
  localparam th_myfunc_42_11 = 11;
  localparam th_myfunc_42_12 = 12;
  localparam th_myfunc_42_13 = 13;
  localparam th_myfunc_42_14 = 14;
  localparam th_myfunc_42_15 = 15;
  localparam th_myfunc_42_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_42 <= th_myfunc_42_init;
      _th_myfunc_42_called <= 0;
      _th_myfunc_42_tid_535 <= 0;
      _th_myfunc_42_tid_536 <= 0;
      _th_myfunc_42_time_537 <= 0;
      _th_myfunc_42_i_538 <= 0;
      _th_myfunc_42___539 <= 0;
    end else begin
      case(th_myfunc_42)
        th_myfunc_42_init: begin
          if(_th_myfunc_start[42] && (th_blink == 10)) begin
            _th_myfunc_42_called <= 1;
          end 
          if(_th_myfunc_start[42] && (th_blink == 10)) begin
            _th_myfunc_42_tid_535 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[42]) begin
            th_myfunc_42 <= th_myfunc_42_1;
          end 
        end
        th_myfunc_42_1: begin
          _th_myfunc_42_tid_536 <= _th_myfunc_42_tid_535;
          th_myfunc_42 <= th_myfunc_42_2;
        end
        th_myfunc_42_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 42)) begin
            th_myfunc_42 <= th_myfunc_42_3;
          end 
        end
        th_myfunc_42_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 42))) begin
            th_myfunc_42 <= th_myfunc_42_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 42)) begin
            th_myfunc_42 <= th_myfunc_42_4;
          end 
        end
        th_myfunc_42_4: begin
          $display("Thread %d Lock", _th_myfunc_42_tid_536);
          th_myfunc_42 <= th_myfunc_42_5;
        end
        th_myfunc_42_5: begin
          _th_myfunc_42_time_537 <= sw;
          th_myfunc_42 <= th_myfunc_42_6;
        end
        th_myfunc_42_6: begin
          _th_myfunc_42_i_538 <= 0;
          th_myfunc_42 <= th_myfunc_42_7;
        end
        th_myfunc_42_7: begin
          if(_th_myfunc_42_i_538 < _th_myfunc_42_time_537) begin
            th_myfunc_42 <= th_myfunc_42_8;
          end else begin
            th_myfunc_42 <= th_myfunc_42_12;
          end
        end
        th_myfunc_42_8: begin
          _th_myfunc_42___539 <= 0;
          th_myfunc_42 <= th_myfunc_42_9;
        end
        th_myfunc_42_9: begin
          if(_th_myfunc_42___539 < 1024) begin
            th_myfunc_42 <= th_myfunc_42_10;
          end else begin
            th_myfunc_42 <= th_myfunc_42_11;
          end
        end
        th_myfunc_42_10: begin
          _th_myfunc_42___539 <= _th_myfunc_42___539 + 1;
          th_myfunc_42 <= th_myfunc_42_9;
        end
        th_myfunc_42_11: begin
          _th_myfunc_42_i_538 <= _th_myfunc_42_i_538 + 1;
          th_myfunc_42 <= th_myfunc_42_7;
        end
        th_myfunc_42_12: begin
          th_myfunc_42 <= th_myfunc_42_13;
        end
        th_myfunc_42_13: begin
          $display("Thread %d count = %d", _th_myfunc_42_tid_536, count);
          th_myfunc_42 <= th_myfunc_42_14;
        end
        th_myfunc_42_14: begin
          th_myfunc_42 <= th_myfunc_42_15;
        end
        th_myfunc_42_15: begin
          $display("Thread %d Unlock", _th_myfunc_42_tid_536);
          th_myfunc_42 <= th_myfunc_42_16;
        end
        th_myfunc_42_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 42)) begin
            _th_myfunc_42_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 42)) begin
            th_myfunc_42 <= th_myfunc_42_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_43_1 = 1;
  localparam th_myfunc_43_2 = 2;
  localparam th_myfunc_43_3 = 3;
  localparam th_myfunc_43_4 = 4;
  localparam th_myfunc_43_5 = 5;
  localparam th_myfunc_43_6 = 6;
  localparam th_myfunc_43_7 = 7;
  localparam th_myfunc_43_8 = 8;
  localparam th_myfunc_43_9 = 9;
  localparam th_myfunc_43_10 = 10;
  localparam th_myfunc_43_11 = 11;
  localparam th_myfunc_43_12 = 12;
  localparam th_myfunc_43_13 = 13;
  localparam th_myfunc_43_14 = 14;
  localparam th_myfunc_43_15 = 15;
  localparam th_myfunc_43_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_43 <= th_myfunc_43_init;
      _th_myfunc_43_called <= 0;
      _th_myfunc_43_tid_540 <= 0;
      _th_myfunc_43_tid_541 <= 0;
      _th_myfunc_43_time_542 <= 0;
      _th_myfunc_43_i_543 <= 0;
      _th_myfunc_43___544 <= 0;
    end else begin
      case(th_myfunc_43)
        th_myfunc_43_init: begin
          if(_th_myfunc_start[43] && (th_blink == 10)) begin
            _th_myfunc_43_called <= 1;
          end 
          if(_th_myfunc_start[43] && (th_blink == 10)) begin
            _th_myfunc_43_tid_540 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[43]) begin
            th_myfunc_43 <= th_myfunc_43_1;
          end 
        end
        th_myfunc_43_1: begin
          _th_myfunc_43_tid_541 <= _th_myfunc_43_tid_540;
          th_myfunc_43 <= th_myfunc_43_2;
        end
        th_myfunc_43_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 43)) begin
            th_myfunc_43 <= th_myfunc_43_3;
          end 
        end
        th_myfunc_43_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 43))) begin
            th_myfunc_43 <= th_myfunc_43_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 43)) begin
            th_myfunc_43 <= th_myfunc_43_4;
          end 
        end
        th_myfunc_43_4: begin
          $display("Thread %d Lock", _th_myfunc_43_tid_541);
          th_myfunc_43 <= th_myfunc_43_5;
        end
        th_myfunc_43_5: begin
          _th_myfunc_43_time_542 <= sw;
          th_myfunc_43 <= th_myfunc_43_6;
        end
        th_myfunc_43_6: begin
          _th_myfunc_43_i_543 <= 0;
          th_myfunc_43 <= th_myfunc_43_7;
        end
        th_myfunc_43_7: begin
          if(_th_myfunc_43_i_543 < _th_myfunc_43_time_542) begin
            th_myfunc_43 <= th_myfunc_43_8;
          end else begin
            th_myfunc_43 <= th_myfunc_43_12;
          end
        end
        th_myfunc_43_8: begin
          _th_myfunc_43___544 <= 0;
          th_myfunc_43 <= th_myfunc_43_9;
        end
        th_myfunc_43_9: begin
          if(_th_myfunc_43___544 < 1024) begin
            th_myfunc_43 <= th_myfunc_43_10;
          end else begin
            th_myfunc_43 <= th_myfunc_43_11;
          end
        end
        th_myfunc_43_10: begin
          _th_myfunc_43___544 <= _th_myfunc_43___544 + 1;
          th_myfunc_43 <= th_myfunc_43_9;
        end
        th_myfunc_43_11: begin
          _th_myfunc_43_i_543 <= _th_myfunc_43_i_543 + 1;
          th_myfunc_43 <= th_myfunc_43_7;
        end
        th_myfunc_43_12: begin
          th_myfunc_43 <= th_myfunc_43_13;
        end
        th_myfunc_43_13: begin
          $display("Thread %d count = %d", _th_myfunc_43_tid_541, count);
          th_myfunc_43 <= th_myfunc_43_14;
        end
        th_myfunc_43_14: begin
          th_myfunc_43 <= th_myfunc_43_15;
        end
        th_myfunc_43_15: begin
          $display("Thread %d Unlock", _th_myfunc_43_tid_541);
          th_myfunc_43 <= th_myfunc_43_16;
        end
        th_myfunc_43_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 43)) begin
            _th_myfunc_43_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 43)) begin
            th_myfunc_43 <= th_myfunc_43_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_44_1 = 1;
  localparam th_myfunc_44_2 = 2;
  localparam th_myfunc_44_3 = 3;
  localparam th_myfunc_44_4 = 4;
  localparam th_myfunc_44_5 = 5;
  localparam th_myfunc_44_6 = 6;
  localparam th_myfunc_44_7 = 7;
  localparam th_myfunc_44_8 = 8;
  localparam th_myfunc_44_9 = 9;
  localparam th_myfunc_44_10 = 10;
  localparam th_myfunc_44_11 = 11;
  localparam th_myfunc_44_12 = 12;
  localparam th_myfunc_44_13 = 13;
  localparam th_myfunc_44_14 = 14;
  localparam th_myfunc_44_15 = 15;
  localparam th_myfunc_44_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_44 <= th_myfunc_44_init;
      _th_myfunc_44_called <= 0;
      _th_myfunc_44_tid_545 <= 0;
      _th_myfunc_44_tid_546 <= 0;
      _th_myfunc_44_time_547 <= 0;
      _th_myfunc_44_i_548 <= 0;
      _th_myfunc_44___549 <= 0;
    end else begin
      case(th_myfunc_44)
        th_myfunc_44_init: begin
          if(_th_myfunc_start[44] && (th_blink == 10)) begin
            _th_myfunc_44_called <= 1;
          end 
          if(_th_myfunc_start[44] && (th_blink == 10)) begin
            _th_myfunc_44_tid_545 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[44]) begin
            th_myfunc_44 <= th_myfunc_44_1;
          end 
        end
        th_myfunc_44_1: begin
          _th_myfunc_44_tid_546 <= _th_myfunc_44_tid_545;
          th_myfunc_44 <= th_myfunc_44_2;
        end
        th_myfunc_44_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 44)) begin
            th_myfunc_44 <= th_myfunc_44_3;
          end 
        end
        th_myfunc_44_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 44))) begin
            th_myfunc_44 <= th_myfunc_44_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 44)) begin
            th_myfunc_44 <= th_myfunc_44_4;
          end 
        end
        th_myfunc_44_4: begin
          $display("Thread %d Lock", _th_myfunc_44_tid_546);
          th_myfunc_44 <= th_myfunc_44_5;
        end
        th_myfunc_44_5: begin
          _th_myfunc_44_time_547 <= sw;
          th_myfunc_44 <= th_myfunc_44_6;
        end
        th_myfunc_44_6: begin
          _th_myfunc_44_i_548 <= 0;
          th_myfunc_44 <= th_myfunc_44_7;
        end
        th_myfunc_44_7: begin
          if(_th_myfunc_44_i_548 < _th_myfunc_44_time_547) begin
            th_myfunc_44 <= th_myfunc_44_8;
          end else begin
            th_myfunc_44 <= th_myfunc_44_12;
          end
        end
        th_myfunc_44_8: begin
          _th_myfunc_44___549 <= 0;
          th_myfunc_44 <= th_myfunc_44_9;
        end
        th_myfunc_44_9: begin
          if(_th_myfunc_44___549 < 1024) begin
            th_myfunc_44 <= th_myfunc_44_10;
          end else begin
            th_myfunc_44 <= th_myfunc_44_11;
          end
        end
        th_myfunc_44_10: begin
          _th_myfunc_44___549 <= _th_myfunc_44___549 + 1;
          th_myfunc_44 <= th_myfunc_44_9;
        end
        th_myfunc_44_11: begin
          _th_myfunc_44_i_548 <= _th_myfunc_44_i_548 + 1;
          th_myfunc_44 <= th_myfunc_44_7;
        end
        th_myfunc_44_12: begin
          th_myfunc_44 <= th_myfunc_44_13;
        end
        th_myfunc_44_13: begin
          $display("Thread %d count = %d", _th_myfunc_44_tid_546, count);
          th_myfunc_44 <= th_myfunc_44_14;
        end
        th_myfunc_44_14: begin
          th_myfunc_44 <= th_myfunc_44_15;
        end
        th_myfunc_44_15: begin
          $display("Thread %d Unlock", _th_myfunc_44_tid_546);
          th_myfunc_44 <= th_myfunc_44_16;
        end
        th_myfunc_44_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 44)) begin
            _th_myfunc_44_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 44)) begin
            th_myfunc_44 <= th_myfunc_44_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_45_1 = 1;
  localparam th_myfunc_45_2 = 2;
  localparam th_myfunc_45_3 = 3;
  localparam th_myfunc_45_4 = 4;
  localparam th_myfunc_45_5 = 5;
  localparam th_myfunc_45_6 = 6;
  localparam th_myfunc_45_7 = 7;
  localparam th_myfunc_45_8 = 8;
  localparam th_myfunc_45_9 = 9;
  localparam th_myfunc_45_10 = 10;
  localparam th_myfunc_45_11 = 11;
  localparam th_myfunc_45_12 = 12;
  localparam th_myfunc_45_13 = 13;
  localparam th_myfunc_45_14 = 14;
  localparam th_myfunc_45_15 = 15;
  localparam th_myfunc_45_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_45 <= th_myfunc_45_init;
      _th_myfunc_45_called <= 0;
      _th_myfunc_45_tid_550 <= 0;
      _th_myfunc_45_tid_551 <= 0;
      _th_myfunc_45_time_552 <= 0;
      _th_myfunc_45_i_553 <= 0;
      _th_myfunc_45___554 <= 0;
    end else begin
      case(th_myfunc_45)
        th_myfunc_45_init: begin
          if(_th_myfunc_start[45] && (th_blink == 10)) begin
            _th_myfunc_45_called <= 1;
          end 
          if(_th_myfunc_start[45] && (th_blink == 10)) begin
            _th_myfunc_45_tid_550 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[45]) begin
            th_myfunc_45 <= th_myfunc_45_1;
          end 
        end
        th_myfunc_45_1: begin
          _th_myfunc_45_tid_551 <= _th_myfunc_45_tid_550;
          th_myfunc_45 <= th_myfunc_45_2;
        end
        th_myfunc_45_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 45)) begin
            th_myfunc_45 <= th_myfunc_45_3;
          end 
        end
        th_myfunc_45_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 45))) begin
            th_myfunc_45 <= th_myfunc_45_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 45)) begin
            th_myfunc_45 <= th_myfunc_45_4;
          end 
        end
        th_myfunc_45_4: begin
          $display("Thread %d Lock", _th_myfunc_45_tid_551);
          th_myfunc_45 <= th_myfunc_45_5;
        end
        th_myfunc_45_5: begin
          _th_myfunc_45_time_552 <= sw;
          th_myfunc_45 <= th_myfunc_45_6;
        end
        th_myfunc_45_6: begin
          _th_myfunc_45_i_553 <= 0;
          th_myfunc_45 <= th_myfunc_45_7;
        end
        th_myfunc_45_7: begin
          if(_th_myfunc_45_i_553 < _th_myfunc_45_time_552) begin
            th_myfunc_45 <= th_myfunc_45_8;
          end else begin
            th_myfunc_45 <= th_myfunc_45_12;
          end
        end
        th_myfunc_45_8: begin
          _th_myfunc_45___554 <= 0;
          th_myfunc_45 <= th_myfunc_45_9;
        end
        th_myfunc_45_9: begin
          if(_th_myfunc_45___554 < 1024) begin
            th_myfunc_45 <= th_myfunc_45_10;
          end else begin
            th_myfunc_45 <= th_myfunc_45_11;
          end
        end
        th_myfunc_45_10: begin
          _th_myfunc_45___554 <= _th_myfunc_45___554 + 1;
          th_myfunc_45 <= th_myfunc_45_9;
        end
        th_myfunc_45_11: begin
          _th_myfunc_45_i_553 <= _th_myfunc_45_i_553 + 1;
          th_myfunc_45 <= th_myfunc_45_7;
        end
        th_myfunc_45_12: begin
          th_myfunc_45 <= th_myfunc_45_13;
        end
        th_myfunc_45_13: begin
          $display("Thread %d count = %d", _th_myfunc_45_tid_551, count);
          th_myfunc_45 <= th_myfunc_45_14;
        end
        th_myfunc_45_14: begin
          th_myfunc_45 <= th_myfunc_45_15;
        end
        th_myfunc_45_15: begin
          $display("Thread %d Unlock", _th_myfunc_45_tid_551);
          th_myfunc_45 <= th_myfunc_45_16;
        end
        th_myfunc_45_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 45)) begin
            _th_myfunc_45_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 45)) begin
            th_myfunc_45 <= th_myfunc_45_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_46_1 = 1;
  localparam th_myfunc_46_2 = 2;
  localparam th_myfunc_46_3 = 3;
  localparam th_myfunc_46_4 = 4;
  localparam th_myfunc_46_5 = 5;
  localparam th_myfunc_46_6 = 6;
  localparam th_myfunc_46_7 = 7;
  localparam th_myfunc_46_8 = 8;
  localparam th_myfunc_46_9 = 9;
  localparam th_myfunc_46_10 = 10;
  localparam th_myfunc_46_11 = 11;
  localparam th_myfunc_46_12 = 12;
  localparam th_myfunc_46_13 = 13;
  localparam th_myfunc_46_14 = 14;
  localparam th_myfunc_46_15 = 15;
  localparam th_myfunc_46_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_46 <= th_myfunc_46_init;
      _th_myfunc_46_called <= 0;
      _th_myfunc_46_tid_555 <= 0;
      _th_myfunc_46_tid_556 <= 0;
      _th_myfunc_46_time_557 <= 0;
      _th_myfunc_46_i_558 <= 0;
      _th_myfunc_46___559 <= 0;
    end else begin
      case(th_myfunc_46)
        th_myfunc_46_init: begin
          if(_th_myfunc_start[46] && (th_blink == 10)) begin
            _th_myfunc_46_called <= 1;
          end 
          if(_th_myfunc_start[46] && (th_blink == 10)) begin
            _th_myfunc_46_tid_555 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[46]) begin
            th_myfunc_46 <= th_myfunc_46_1;
          end 
        end
        th_myfunc_46_1: begin
          _th_myfunc_46_tid_556 <= _th_myfunc_46_tid_555;
          th_myfunc_46 <= th_myfunc_46_2;
        end
        th_myfunc_46_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 46)) begin
            th_myfunc_46 <= th_myfunc_46_3;
          end 
        end
        th_myfunc_46_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 46))) begin
            th_myfunc_46 <= th_myfunc_46_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 46)) begin
            th_myfunc_46 <= th_myfunc_46_4;
          end 
        end
        th_myfunc_46_4: begin
          $display("Thread %d Lock", _th_myfunc_46_tid_556);
          th_myfunc_46 <= th_myfunc_46_5;
        end
        th_myfunc_46_5: begin
          _th_myfunc_46_time_557 <= sw;
          th_myfunc_46 <= th_myfunc_46_6;
        end
        th_myfunc_46_6: begin
          _th_myfunc_46_i_558 <= 0;
          th_myfunc_46 <= th_myfunc_46_7;
        end
        th_myfunc_46_7: begin
          if(_th_myfunc_46_i_558 < _th_myfunc_46_time_557) begin
            th_myfunc_46 <= th_myfunc_46_8;
          end else begin
            th_myfunc_46 <= th_myfunc_46_12;
          end
        end
        th_myfunc_46_8: begin
          _th_myfunc_46___559 <= 0;
          th_myfunc_46 <= th_myfunc_46_9;
        end
        th_myfunc_46_9: begin
          if(_th_myfunc_46___559 < 1024) begin
            th_myfunc_46 <= th_myfunc_46_10;
          end else begin
            th_myfunc_46 <= th_myfunc_46_11;
          end
        end
        th_myfunc_46_10: begin
          _th_myfunc_46___559 <= _th_myfunc_46___559 + 1;
          th_myfunc_46 <= th_myfunc_46_9;
        end
        th_myfunc_46_11: begin
          _th_myfunc_46_i_558 <= _th_myfunc_46_i_558 + 1;
          th_myfunc_46 <= th_myfunc_46_7;
        end
        th_myfunc_46_12: begin
          th_myfunc_46 <= th_myfunc_46_13;
        end
        th_myfunc_46_13: begin
          $display("Thread %d count = %d", _th_myfunc_46_tid_556, count);
          th_myfunc_46 <= th_myfunc_46_14;
        end
        th_myfunc_46_14: begin
          th_myfunc_46 <= th_myfunc_46_15;
        end
        th_myfunc_46_15: begin
          $display("Thread %d Unlock", _th_myfunc_46_tid_556);
          th_myfunc_46 <= th_myfunc_46_16;
        end
        th_myfunc_46_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 46)) begin
            _th_myfunc_46_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 46)) begin
            th_myfunc_46 <= th_myfunc_46_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_47_1 = 1;
  localparam th_myfunc_47_2 = 2;
  localparam th_myfunc_47_3 = 3;
  localparam th_myfunc_47_4 = 4;
  localparam th_myfunc_47_5 = 5;
  localparam th_myfunc_47_6 = 6;
  localparam th_myfunc_47_7 = 7;
  localparam th_myfunc_47_8 = 8;
  localparam th_myfunc_47_9 = 9;
  localparam th_myfunc_47_10 = 10;
  localparam th_myfunc_47_11 = 11;
  localparam th_myfunc_47_12 = 12;
  localparam th_myfunc_47_13 = 13;
  localparam th_myfunc_47_14 = 14;
  localparam th_myfunc_47_15 = 15;
  localparam th_myfunc_47_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_47 <= th_myfunc_47_init;
      _th_myfunc_47_called <= 0;
      _th_myfunc_47_tid_560 <= 0;
      _th_myfunc_47_tid_561 <= 0;
      _th_myfunc_47_time_562 <= 0;
      _th_myfunc_47_i_563 <= 0;
      _th_myfunc_47___564 <= 0;
    end else begin
      case(th_myfunc_47)
        th_myfunc_47_init: begin
          if(_th_myfunc_start[47] && (th_blink == 10)) begin
            _th_myfunc_47_called <= 1;
          end 
          if(_th_myfunc_start[47] && (th_blink == 10)) begin
            _th_myfunc_47_tid_560 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[47]) begin
            th_myfunc_47 <= th_myfunc_47_1;
          end 
        end
        th_myfunc_47_1: begin
          _th_myfunc_47_tid_561 <= _th_myfunc_47_tid_560;
          th_myfunc_47 <= th_myfunc_47_2;
        end
        th_myfunc_47_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 47)) begin
            th_myfunc_47 <= th_myfunc_47_3;
          end 
        end
        th_myfunc_47_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 47))) begin
            th_myfunc_47 <= th_myfunc_47_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 47)) begin
            th_myfunc_47 <= th_myfunc_47_4;
          end 
        end
        th_myfunc_47_4: begin
          $display("Thread %d Lock", _th_myfunc_47_tid_561);
          th_myfunc_47 <= th_myfunc_47_5;
        end
        th_myfunc_47_5: begin
          _th_myfunc_47_time_562 <= sw;
          th_myfunc_47 <= th_myfunc_47_6;
        end
        th_myfunc_47_6: begin
          _th_myfunc_47_i_563 <= 0;
          th_myfunc_47 <= th_myfunc_47_7;
        end
        th_myfunc_47_7: begin
          if(_th_myfunc_47_i_563 < _th_myfunc_47_time_562) begin
            th_myfunc_47 <= th_myfunc_47_8;
          end else begin
            th_myfunc_47 <= th_myfunc_47_12;
          end
        end
        th_myfunc_47_8: begin
          _th_myfunc_47___564 <= 0;
          th_myfunc_47 <= th_myfunc_47_9;
        end
        th_myfunc_47_9: begin
          if(_th_myfunc_47___564 < 1024) begin
            th_myfunc_47 <= th_myfunc_47_10;
          end else begin
            th_myfunc_47 <= th_myfunc_47_11;
          end
        end
        th_myfunc_47_10: begin
          _th_myfunc_47___564 <= _th_myfunc_47___564 + 1;
          th_myfunc_47 <= th_myfunc_47_9;
        end
        th_myfunc_47_11: begin
          _th_myfunc_47_i_563 <= _th_myfunc_47_i_563 + 1;
          th_myfunc_47 <= th_myfunc_47_7;
        end
        th_myfunc_47_12: begin
          th_myfunc_47 <= th_myfunc_47_13;
        end
        th_myfunc_47_13: begin
          $display("Thread %d count = %d", _th_myfunc_47_tid_561, count);
          th_myfunc_47 <= th_myfunc_47_14;
        end
        th_myfunc_47_14: begin
          th_myfunc_47 <= th_myfunc_47_15;
        end
        th_myfunc_47_15: begin
          $display("Thread %d Unlock", _th_myfunc_47_tid_561);
          th_myfunc_47 <= th_myfunc_47_16;
        end
        th_myfunc_47_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 47)) begin
            _th_myfunc_47_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 47)) begin
            th_myfunc_47 <= th_myfunc_47_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_48_1 = 1;
  localparam th_myfunc_48_2 = 2;
  localparam th_myfunc_48_3 = 3;
  localparam th_myfunc_48_4 = 4;
  localparam th_myfunc_48_5 = 5;
  localparam th_myfunc_48_6 = 6;
  localparam th_myfunc_48_7 = 7;
  localparam th_myfunc_48_8 = 8;
  localparam th_myfunc_48_9 = 9;
  localparam th_myfunc_48_10 = 10;
  localparam th_myfunc_48_11 = 11;
  localparam th_myfunc_48_12 = 12;
  localparam th_myfunc_48_13 = 13;
  localparam th_myfunc_48_14 = 14;
  localparam th_myfunc_48_15 = 15;
  localparam th_myfunc_48_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_48 <= th_myfunc_48_init;
      _th_myfunc_48_called <= 0;
      _th_myfunc_48_tid_565 <= 0;
      _th_myfunc_48_tid_566 <= 0;
      _th_myfunc_48_time_567 <= 0;
      _th_myfunc_48_i_568 <= 0;
      _th_myfunc_48___569 <= 0;
    end else begin
      case(th_myfunc_48)
        th_myfunc_48_init: begin
          if(_th_myfunc_start[48] && (th_blink == 10)) begin
            _th_myfunc_48_called <= 1;
          end 
          if(_th_myfunc_start[48] && (th_blink == 10)) begin
            _th_myfunc_48_tid_565 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[48]) begin
            th_myfunc_48 <= th_myfunc_48_1;
          end 
        end
        th_myfunc_48_1: begin
          _th_myfunc_48_tid_566 <= _th_myfunc_48_tid_565;
          th_myfunc_48 <= th_myfunc_48_2;
        end
        th_myfunc_48_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 48)) begin
            th_myfunc_48 <= th_myfunc_48_3;
          end 
        end
        th_myfunc_48_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 48))) begin
            th_myfunc_48 <= th_myfunc_48_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 48)) begin
            th_myfunc_48 <= th_myfunc_48_4;
          end 
        end
        th_myfunc_48_4: begin
          $display("Thread %d Lock", _th_myfunc_48_tid_566);
          th_myfunc_48 <= th_myfunc_48_5;
        end
        th_myfunc_48_5: begin
          _th_myfunc_48_time_567 <= sw;
          th_myfunc_48 <= th_myfunc_48_6;
        end
        th_myfunc_48_6: begin
          _th_myfunc_48_i_568 <= 0;
          th_myfunc_48 <= th_myfunc_48_7;
        end
        th_myfunc_48_7: begin
          if(_th_myfunc_48_i_568 < _th_myfunc_48_time_567) begin
            th_myfunc_48 <= th_myfunc_48_8;
          end else begin
            th_myfunc_48 <= th_myfunc_48_12;
          end
        end
        th_myfunc_48_8: begin
          _th_myfunc_48___569 <= 0;
          th_myfunc_48 <= th_myfunc_48_9;
        end
        th_myfunc_48_9: begin
          if(_th_myfunc_48___569 < 1024) begin
            th_myfunc_48 <= th_myfunc_48_10;
          end else begin
            th_myfunc_48 <= th_myfunc_48_11;
          end
        end
        th_myfunc_48_10: begin
          _th_myfunc_48___569 <= _th_myfunc_48___569 + 1;
          th_myfunc_48 <= th_myfunc_48_9;
        end
        th_myfunc_48_11: begin
          _th_myfunc_48_i_568 <= _th_myfunc_48_i_568 + 1;
          th_myfunc_48 <= th_myfunc_48_7;
        end
        th_myfunc_48_12: begin
          th_myfunc_48 <= th_myfunc_48_13;
        end
        th_myfunc_48_13: begin
          $display("Thread %d count = %d", _th_myfunc_48_tid_566, count);
          th_myfunc_48 <= th_myfunc_48_14;
        end
        th_myfunc_48_14: begin
          th_myfunc_48 <= th_myfunc_48_15;
        end
        th_myfunc_48_15: begin
          $display("Thread %d Unlock", _th_myfunc_48_tid_566);
          th_myfunc_48 <= th_myfunc_48_16;
        end
        th_myfunc_48_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 48)) begin
            _th_myfunc_48_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 48)) begin
            th_myfunc_48 <= th_myfunc_48_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_49_1 = 1;
  localparam th_myfunc_49_2 = 2;
  localparam th_myfunc_49_3 = 3;
  localparam th_myfunc_49_4 = 4;
  localparam th_myfunc_49_5 = 5;
  localparam th_myfunc_49_6 = 6;
  localparam th_myfunc_49_7 = 7;
  localparam th_myfunc_49_8 = 8;
  localparam th_myfunc_49_9 = 9;
  localparam th_myfunc_49_10 = 10;
  localparam th_myfunc_49_11 = 11;
  localparam th_myfunc_49_12 = 12;
  localparam th_myfunc_49_13 = 13;
  localparam th_myfunc_49_14 = 14;
  localparam th_myfunc_49_15 = 15;
  localparam th_myfunc_49_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_49 <= th_myfunc_49_init;
      _th_myfunc_49_called <= 0;
      _th_myfunc_49_tid_570 <= 0;
      _th_myfunc_49_tid_571 <= 0;
      _th_myfunc_49_time_572 <= 0;
      _th_myfunc_49_i_573 <= 0;
      _th_myfunc_49___574 <= 0;
    end else begin
      case(th_myfunc_49)
        th_myfunc_49_init: begin
          if(_th_myfunc_start[49] && (th_blink == 10)) begin
            _th_myfunc_49_called <= 1;
          end 
          if(_th_myfunc_start[49] && (th_blink == 10)) begin
            _th_myfunc_49_tid_570 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[49]) begin
            th_myfunc_49 <= th_myfunc_49_1;
          end 
        end
        th_myfunc_49_1: begin
          _th_myfunc_49_tid_571 <= _th_myfunc_49_tid_570;
          th_myfunc_49 <= th_myfunc_49_2;
        end
        th_myfunc_49_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 49)) begin
            th_myfunc_49 <= th_myfunc_49_3;
          end 
        end
        th_myfunc_49_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 49))) begin
            th_myfunc_49 <= th_myfunc_49_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 49)) begin
            th_myfunc_49 <= th_myfunc_49_4;
          end 
        end
        th_myfunc_49_4: begin
          $display("Thread %d Lock", _th_myfunc_49_tid_571);
          th_myfunc_49 <= th_myfunc_49_5;
        end
        th_myfunc_49_5: begin
          _th_myfunc_49_time_572 <= sw;
          th_myfunc_49 <= th_myfunc_49_6;
        end
        th_myfunc_49_6: begin
          _th_myfunc_49_i_573 <= 0;
          th_myfunc_49 <= th_myfunc_49_7;
        end
        th_myfunc_49_7: begin
          if(_th_myfunc_49_i_573 < _th_myfunc_49_time_572) begin
            th_myfunc_49 <= th_myfunc_49_8;
          end else begin
            th_myfunc_49 <= th_myfunc_49_12;
          end
        end
        th_myfunc_49_8: begin
          _th_myfunc_49___574 <= 0;
          th_myfunc_49 <= th_myfunc_49_9;
        end
        th_myfunc_49_9: begin
          if(_th_myfunc_49___574 < 1024) begin
            th_myfunc_49 <= th_myfunc_49_10;
          end else begin
            th_myfunc_49 <= th_myfunc_49_11;
          end
        end
        th_myfunc_49_10: begin
          _th_myfunc_49___574 <= _th_myfunc_49___574 + 1;
          th_myfunc_49 <= th_myfunc_49_9;
        end
        th_myfunc_49_11: begin
          _th_myfunc_49_i_573 <= _th_myfunc_49_i_573 + 1;
          th_myfunc_49 <= th_myfunc_49_7;
        end
        th_myfunc_49_12: begin
          th_myfunc_49 <= th_myfunc_49_13;
        end
        th_myfunc_49_13: begin
          $display("Thread %d count = %d", _th_myfunc_49_tid_571, count);
          th_myfunc_49 <= th_myfunc_49_14;
        end
        th_myfunc_49_14: begin
          th_myfunc_49 <= th_myfunc_49_15;
        end
        th_myfunc_49_15: begin
          $display("Thread %d Unlock", _th_myfunc_49_tid_571);
          th_myfunc_49 <= th_myfunc_49_16;
        end
        th_myfunc_49_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 49)) begin
            _th_myfunc_49_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 49)) begin
            th_myfunc_49 <= th_myfunc_49_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_50_1 = 1;
  localparam th_myfunc_50_2 = 2;
  localparam th_myfunc_50_3 = 3;
  localparam th_myfunc_50_4 = 4;
  localparam th_myfunc_50_5 = 5;
  localparam th_myfunc_50_6 = 6;
  localparam th_myfunc_50_7 = 7;
  localparam th_myfunc_50_8 = 8;
  localparam th_myfunc_50_9 = 9;
  localparam th_myfunc_50_10 = 10;
  localparam th_myfunc_50_11 = 11;
  localparam th_myfunc_50_12 = 12;
  localparam th_myfunc_50_13 = 13;
  localparam th_myfunc_50_14 = 14;
  localparam th_myfunc_50_15 = 15;
  localparam th_myfunc_50_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_50 <= th_myfunc_50_init;
      _th_myfunc_50_called <= 0;
      _th_myfunc_50_tid_575 <= 0;
      _th_myfunc_50_tid_576 <= 0;
      _th_myfunc_50_time_577 <= 0;
      _th_myfunc_50_i_578 <= 0;
      _th_myfunc_50___579 <= 0;
    end else begin
      case(th_myfunc_50)
        th_myfunc_50_init: begin
          if(_th_myfunc_start[50] && (th_blink == 10)) begin
            _th_myfunc_50_called <= 1;
          end 
          if(_th_myfunc_start[50] && (th_blink == 10)) begin
            _th_myfunc_50_tid_575 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[50]) begin
            th_myfunc_50 <= th_myfunc_50_1;
          end 
        end
        th_myfunc_50_1: begin
          _th_myfunc_50_tid_576 <= _th_myfunc_50_tid_575;
          th_myfunc_50 <= th_myfunc_50_2;
        end
        th_myfunc_50_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 50)) begin
            th_myfunc_50 <= th_myfunc_50_3;
          end 
        end
        th_myfunc_50_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 50))) begin
            th_myfunc_50 <= th_myfunc_50_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 50)) begin
            th_myfunc_50 <= th_myfunc_50_4;
          end 
        end
        th_myfunc_50_4: begin
          $display("Thread %d Lock", _th_myfunc_50_tid_576);
          th_myfunc_50 <= th_myfunc_50_5;
        end
        th_myfunc_50_5: begin
          _th_myfunc_50_time_577 <= sw;
          th_myfunc_50 <= th_myfunc_50_6;
        end
        th_myfunc_50_6: begin
          _th_myfunc_50_i_578 <= 0;
          th_myfunc_50 <= th_myfunc_50_7;
        end
        th_myfunc_50_7: begin
          if(_th_myfunc_50_i_578 < _th_myfunc_50_time_577) begin
            th_myfunc_50 <= th_myfunc_50_8;
          end else begin
            th_myfunc_50 <= th_myfunc_50_12;
          end
        end
        th_myfunc_50_8: begin
          _th_myfunc_50___579 <= 0;
          th_myfunc_50 <= th_myfunc_50_9;
        end
        th_myfunc_50_9: begin
          if(_th_myfunc_50___579 < 1024) begin
            th_myfunc_50 <= th_myfunc_50_10;
          end else begin
            th_myfunc_50 <= th_myfunc_50_11;
          end
        end
        th_myfunc_50_10: begin
          _th_myfunc_50___579 <= _th_myfunc_50___579 + 1;
          th_myfunc_50 <= th_myfunc_50_9;
        end
        th_myfunc_50_11: begin
          _th_myfunc_50_i_578 <= _th_myfunc_50_i_578 + 1;
          th_myfunc_50 <= th_myfunc_50_7;
        end
        th_myfunc_50_12: begin
          th_myfunc_50 <= th_myfunc_50_13;
        end
        th_myfunc_50_13: begin
          $display("Thread %d count = %d", _th_myfunc_50_tid_576, count);
          th_myfunc_50 <= th_myfunc_50_14;
        end
        th_myfunc_50_14: begin
          th_myfunc_50 <= th_myfunc_50_15;
        end
        th_myfunc_50_15: begin
          $display("Thread %d Unlock", _th_myfunc_50_tid_576);
          th_myfunc_50 <= th_myfunc_50_16;
        end
        th_myfunc_50_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 50)) begin
            _th_myfunc_50_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 50)) begin
            th_myfunc_50 <= th_myfunc_50_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_51_1 = 1;
  localparam th_myfunc_51_2 = 2;
  localparam th_myfunc_51_3 = 3;
  localparam th_myfunc_51_4 = 4;
  localparam th_myfunc_51_5 = 5;
  localparam th_myfunc_51_6 = 6;
  localparam th_myfunc_51_7 = 7;
  localparam th_myfunc_51_8 = 8;
  localparam th_myfunc_51_9 = 9;
  localparam th_myfunc_51_10 = 10;
  localparam th_myfunc_51_11 = 11;
  localparam th_myfunc_51_12 = 12;
  localparam th_myfunc_51_13 = 13;
  localparam th_myfunc_51_14 = 14;
  localparam th_myfunc_51_15 = 15;
  localparam th_myfunc_51_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_51 <= th_myfunc_51_init;
      _th_myfunc_51_called <= 0;
      _th_myfunc_51_tid_580 <= 0;
      _th_myfunc_51_tid_581 <= 0;
      _th_myfunc_51_time_582 <= 0;
      _th_myfunc_51_i_583 <= 0;
      _th_myfunc_51___584 <= 0;
    end else begin
      case(th_myfunc_51)
        th_myfunc_51_init: begin
          if(_th_myfunc_start[51] && (th_blink == 10)) begin
            _th_myfunc_51_called <= 1;
          end 
          if(_th_myfunc_start[51] && (th_blink == 10)) begin
            _th_myfunc_51_tid_580 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[51]) begin
            th_myfunc_51 <= th_myfunc_51_1;
          end 
        end
        th_myfunc_51_1: begin
          _th_myfunc_51_tid_581 <= _th_myfunc_51_tid_580;
          th_myfunc_51 <= th_myfunc_51_2;
        end
        th_myfunc_51_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 51)) begin
            th_myfunc_51 <= th_myfunc_51_3;
          end 
        end
        th_myfunc_51_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 51))) begin
            th_myfunc_51 <= th_myfunc_51_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 51)) begin
            th_myfunc_51 <= th_myfunc_51_4;
          end 
        end
        th_myfunc_51_4: begin
          $display("Thread %d Lock", _th_myfunc_51_tid_581);
          th_myfunc_51 <= th_myfunc_51_5;
        end
        th_myfunc_51_5: begin
          _th_myfunc_51_time_582 <= sw;
          th_myfunc_51 <= th_myfunc_51_6;
        end
        th_myfunc_51_6: begin
          _th_myfunc_51_i_583 <= 0;
          th_myfunc_51 <= th_myfunc_51_7;
        end
        th_myfunc_51_7: begin
          if(_th_myfunc_51_i_583 < _th_myfunc_51_time_582) begin
            th_myfunc_51 <= th_myfunc_51_8;
          end else begin
            th_myfunc_51 <= th_myfunc_51_12;
          end
        end
        th_myfunc_51_8: begin
          _th_myfunc_51___584 <= 0;
          th_myfunc_51 <= th_myfunc_51_9;
        end
        th_myfunc_51_9: begin
          if(_th_myfunc_51___584 < 1024) begin
            th_myfunc_51 <= th_myfunc_51_10;
          end else begin
            th_myfunc_51 <= th_myfunc_51_11;
          end
        end
        th_myfunc_51_10: begin
          _th_myfunc_51___584 <= _th_myfunc_51___584 + 1;
          th_myfunc_51 <= th_myfunc_51_9;
        end
        th_myfunc_51_11: begin
          _th_myfunc_51_i_583 <= _th_myfunc_51_i_583 + 1;
          th_myfunc_51 <= th_myfunc_51_7;
        end
        th_myfunc_51_12: begin
          th_myfunc_51 <= th_myfunc_51_13;
        end
        th_myfunc_51_13: begin
          $display("Thread %d count = %d", _th_myfunc_51_tid_581, count);
          th_myfunc_51 <= th_myfunc_51_14;
        end
        th_myfunc_51_14: begin
          th_myfunc_51 <= th_myfunc_51_15;
        end
        th_myfunc_51_15: begin
          $display("Thread %d Unlock", _th_myfunc_51_tid_581);
          th_myfunc_51 <= th_myfunc_51_16;
        end
        th_myfunc_51_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 51)) begin
            _th_myfunc_51_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 51)) begin
            th_myfunc_51 <= th_myfunc_51_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_52_1 = 1;
  localparam th_myfunc_52_2 = 2;
  localparam th_myfunc_52_3 = 3;
  localparam th_myfunc_52_4 = 4;
  localparam th_myfunc_52_5 = 5;
  localparam th_myfunc_52_6 = 6;
  localparam th_myfunc_52_7 = 7;
  localparam th_myfunc_52_8 = 8;
  localparam th_myfunc_52_9 = 9;
  localparam th_myfunc_52_10 = 10;
  localparam th_myfunc_52_11 = 11;
  localparam th_myfunc_52_12 = 12;
  localparam th_myfunc_52_13 = 13;
  localparam th_myfunc_52_14 = 14;
  localparam th_myfunc_52_15 = 15;
  localparam th_myfunc_52_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_52 <= th_myfunc_52_init;
      _th_myfunc_52_called <= 0;
      _th_myfunc_52_tid_585 <= 0;
      _th_myfunc_52_tid_586 <= 0;
      _th_myfunc_52_time_587 <= 0;
      _th_myfunc_52_i_588 <= 0;
      _th_myfunc_52___589 <= 0;
    end else begin
      case(th_myfunc_52)
        th_myfunc_52_init: begin
          if(_th_myfunc_start[52] && (th_blink == 10)) begin
            _th_myfunc_52_called <= 1;
          end 
          if(_th_myfunc_start[52] && (th_blink == 10)) begin
            _th_myfunc_52_tid_585 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[52]) begin
            th_myfunc_52 <= th_myfunc_52_1;
          end 
        end
        th_myfunc_52_1: begin
          _th_myfunc_52_tid_586 <= _th_myfunc_52_tid_585;
          th_myfunc_52 <= th_myfunc_52_2;
        end
        th_myfunc_52_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 52)) begin
            th_myfunc_52 <= th_myfunc_52_3;
          end 
        end
        th_myfunc_52_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 52))) begin
            th_myfunc_52 <= th_myfunc_52_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 52)) begin
            th_myfunc_52 <= th_myfunc_52_4;
          end 
        end
        th_myfunc_52_4: begin
          $display("Thread %d Lock", _th_myfunc_52_tid_586);
          th_myfunc_52 <= th_myfunc_52_5;
        end
        th_myfunc_52_5: begin
          _th_myfunc_52_time_587 <= sw;
          th_myfunc_52 <= th_myfunc_52_6;
        end
        th_myfunc_52_6: begin
          _th_myfunc_52_i_588 <= 0;
          th_myfunc_52 <= th_myfunc_52_7;
        end
        th_myfunc_52_7: begin
          if(_th_myfunc_52_i_588 < _th_myfunc_52_time_587) begin
            th_myfunc_52 <= th_myfunc_52_8;
          end else begin
            th_myfunc_52 <= th_myfunc_52_12;
          end
        end
        th_myfunc_52_8: begin
          _th_myfunc_52___589 <= 0;
          th_myfunc_52 <= th_myfunc_52_9;
        end
        th_myfunc_52_9: begin
          if(_th_myfunc_52___589 < 1024) begin
            th_myfunc_52 <= th_myfunc_52_10;
          end else begin
            th_myfunc_52 <= th_myfunc_52_11;
          end
        end
        th_myfunc_52_10: begin
          _th_myfunc_52___589 <= _th_myfunc_52___589 + 1;
          th_myfunc_52 <= th_myfunc_52_9;
        end
        th_myfunc_52_11: begin
          _th_myfunc_52_i_588 <= _th_myfunc_52_i_588 + 1;
          th_myfunc_52 <= th_myfunc_52_7;
        end
        th_myfunc_52_12: begin
          th_myfunc_52 <= th_myfunc_52_13;
        end
        th_myfunc_52_13: begin
          $display("Thread %d count = %d", _th_myfunc_52_tid_586, count);
          th_myfunc_52 <= th_myfunc_52_14;
        end
        th_myfunc_52_14: begin
          th_myfunc_52 <= th_myfunc_52_15;
        end
        th_myfunc_52_15: begin
          $display("Thread %d Unlock", _th_myfunc_52_tid_586);
          th_myfunc_52 <= th_myfunc_52_16;
        end
        th_myfunc_52_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 52)) begin
            _th_myfunc_52_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 52)) begin
            th_myfunc_52 <= th_myfunc_52_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_53_1 = 1;
  localparam th_myfunc_53_2 = 2;
  localparam th_myfunc_53_3 = 3;
  localparam th_myfunc_53_4 = 4;
  localparam th_myfunc_53_5 = 5;
  localparam th_myfunc_53_6 = 6;
  localparam th_myfunc_53_7 = 7;
  localparam th_myfunc_53_8 = 8;
  localparam th_myfunc_53_9 = 9;
  localparam th_myfunc_53_10 = 10;
  localparam th_myfunc_53_11 = 11;
  localparam th_myfunc_53_12 = 12;
  localparam th_myfunc_53_13 = 13;
  localparam th_myfunc_53_14 = 14;
  localparam th_myfunc_53_15 = 15;
  localparam th_myfunc_53_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_53 <= th_myfunc_53_init;
      _th_myfunc_53_called <= 0;
      _th_myfunc_53_tid_590 <= 0;
      _th_myfunc_53_tid_591 <= 0;
      _th_myfunc_53_time_592 <= 0;
      _th_myfunc_53_i_593 <= 0;
      _th_myfunc_53___594 <= 0;
    end else begin
      case(th_myfunc_53)
        th_myfunc_53_init: begin
          if(_th_myfunc_start[53] && (th_blink == 10)) begin
            _th_myfunc_53_called <= 1;
          end 
          if(_th_myfunc_start[53] && (th_blink == 10)) begin
            _th_myfunc_53_tid_590 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[53]) begin
            th_myfunc_53 <= th_myfunc_53_1;
          end 
        end
        th_myfunc_53_1: begin
          _th_myfunc_53_tid_591 <= _th_myfunc_53_tid_590;
          th_myfunc_53 <= th_myfunc_53_2;
        end
        th_myfunc_53_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 53)) begin
            th_myfunc_53 <= th_myfunc_53_3;
          end 
        end
        th_myfunc_53_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 53))) begin
            th_myfunc_53 <= th_myfunc_53_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 53)) begin
            th_myfunc_53 <= th_myfunc_53_4;
          end 
        end
        th_myfunc_53_4: begin
          $display("Thread %d Lock", _th_myfunc_53_tid_591);
          th_myfunc_53 <= th_myfunc_53_5;
        end
        th_myfunc_53_5: begin
          _th_myfunc_53_time_592 <= sw;
          th_myfunc_53 <= th_myfunc_53_6;
        end
        th_myfunc_53_6: begin
          _th_myfunc_53_i_593 <= 0;
          th_myfunc_53 <= th_myfunc_53_7;
        end
        th_myfunc_53_7: begin
          if(_th_myfunc_53_i_593 < _th_myfunc_53_time_592) begin
            th_myfunc_53 <= th_myfunc_53_8;
          end else begin
            th_myfunc_53 <= th_myfunc_53_12;
          end
        end
        th_myfunc_53_8: begin
          _th_myfunc_53___594 <= 0;
          th_myfunc_53 <= th_myfunc_53_9;
        end
        th_myfunc_53_9: begin
          if(_th_myfunc_53___594 < 1024) begin
            th_myfunc_53 <= th_myfunc_53_10;
          end else begin
            th_myfunc_53 <= th_myfunc_53_11;
          end
        end
        th_myfunc_53_10: begin
          _th_myfunc_53___594 <= _th_myfunc_53___594 + 1;
          th_myfunc_53 <= th_myfunc_53_9;
        end
        th_myfunc_53_11: begin
          _th_myfunc_53_i_593 <= _th_myfunc_53_i_593 + 1;
          th_myfunc_53 <= th_myfunc_53_7;
        end
        th_myfunc_53_12: begin
          th_myfunc_53 <= th_myfunc_53_13;
        end
        th_myfunc_53_13: begin
          $display("Thread %d count = %d", _th_myfunc_53_tid_591, count);
          th_myfunc_53 <= th_myfunc_53_14;
        end
        th_myfunc_53_14: begin
          th_myfunc_53 <= th_myfunc_53_15;
        end
        th_myfunc_53_15: begin
          $display("Thread %d Unlock", _th_myfunc_53_tid_591);
          th_myfunc_53 <= th_myfunc_53_16;
        end
        th_myfunc_53_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 53)) begin
            _th_myfunc_53_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 53)) begin
            th_myfunc_53 <= th_myfunc_53_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_54_1 = 1;
  localparam th_myfunc_54_2 = 2;
  localparam th_myfunc_54_3 = 3;
  localparam th_myfunc_54_4 = 4;
  localparam th_myfunc_54_5 = 5;
  localparam th_myfunc_54_6 = 6;
  localparam th_myfunc_54_7 = 7;
  localparam th_myfunc_54_8 = 8;
  localparam th_myfunc_54_9 = 9;
  localparam th_myfunc_54_10 = 10;
  localparam th_myfunc_54_11 = 11;
  localparam th_myfunc_54_12 = 12;
  localparam th_myfunc_54_13 = 13;
  localparam th_myfunc_54_14 = 14;
  localparam th_myfunc_54_15 = 15;
  localparam th_myfunc_54_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_54 <= th_myfunc_54_init;
      _th_myfunc_54_called <= 0;
      _th_myfunc_54_tid_595 <= 0;
      _th_myfunc_54_tid_596 <= 0;
      _th_myfunc_54_time_597 <= 0;
      _th_myfunc_54_i_598 <= 0;
      _th_myfunc_54___599 <= 0;
    end else begin
      case(th_myfunc_54)
        th_myfunc_54_init: begin
          if(_th_myfunc_start[54] && (th_blink == 10)) begin
            _th_myfunc_54_called <= 1;
          end 
          if(_th_myfunc_start[54] && (th_blink == 10)) begin
            _th_myfunc_54_tid_595 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[54]) begin
            th_myfunc_54 <= th_myfunc_54_1;
          end 
        end
        th_myfunc_54_1: begin
          _th_myfunc_54_tid_596 <= _th_myfunc_54_tid_595;
          th_myfunc_54 <= th_myfunc_54_2;
        end
        th_myfunc_54_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 54)) begin
            th_myfunc_54 <= th_myfunc_54_3;
          end 
        end
        th_myfunc_54_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 54))) begin
            th_myfunc_54 <= th_myfunc_54_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 54)) begin
            th_myfunc_54 <= th_myfunc_54_4;
          end 
        end
        th_myfunc_54_4: begin
          $display("Thread %d Lock", _th_myfunc_54_tid_596);
          th_myfunc_54 <= th_myfunc_54_5;
        end
        th_myfunc_54_5: begin
          _th_myfunc_54_time_597 <= sw;
          th_myfunc_54 <= th_myfunc_54_6;
        end
        th_myfunc_54_6: begin
          _th_myfunc_54_i_598 <= 0;
          th_myfunc_54 <= th_myfunc_54_7;
        end
        th_myfunc_54_7: begin
          if(_th_myfunc_54_i_598 < _th_myfunc_54_time_597) begin
            th_myfunc_54 <= th_myfunc_54_8;
          end else begin
            th_myfunc_54 <= th_myfunc_54_12;
          end
        end
        th_myfunc_54_8: begin
          _th_myfunc_54___599 <= 0;
          th_myfunc_54 <= th_myfunc_54_9;
        end
        th_myfunc_54_9: begin
          if(_th_myfunc_54___599 < 1024) begin
            th_myfunc_54 <= th_myfunc_54_10;
          end else begin
            th_myfunc_54 <= th_myfunc_54_11;
          end
        end
        th_myfunc_54_10: begin
          _th_myfunc_54___599 <= _th_myfunc_54___599 + 1;
          th_myfunc_54 <= th_myfunc_54_9;
        end
        th_myfunc_54_11: begin
          _th_myfunc_54_i_598 <= _th_myfunc_54_i_598 + 1;
          th_myfunc_54 <= th_myfunc_54_7;
        end
        th_myfunc_54_12: begin
          th_myfunc_54 <= th_myfunc_54_13;
        end
        th_myfunc_54_13: begin
          $display("Thread %d count = %d", _th_myfunc_54_tid_596, count);
          th_myfunc_54 <= th_myfunc_54_14;
        end
        th_myfunc_54_14: begin
          th_myfunc_54 <= th_myfunc_54_15;
        end
        th_myfunc_54_15: begin
          $display("Thread %d Unlock", _th_myfunc_54_tid_596);
          th_myfunc_54 <= th_myfunc_54_16;
        end
        th_myfunc_54_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 54)) begin
            _th_myfunc_54_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 54)) begin
            th_myfunc_54 <= th_myfunc_54_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_55_1 = 1;
  localparam th_myfunc_55_2 = 2;
  localparam th_myfunc_55_3 = 3;
  localparam th_myfunc_55_4 = 4;
  localparam th_myfunc_55_5 = 5;
  localparam th_myfunc_55_6 = 6;
  localparam th_myfunc_55_7 = 7;
  localparam th_myfunc_55_8 = 8;
  localparam th_myfunc_55_9 = 9;
  localparam th_myfunc_55_10 = 10;
  localparam th_myfunc_55_11 = 11;
  localparam th_myfunc_55_12 = 12;
  localparam th_myfunc_55_13 = 13;
  localparam th_myfunc_55_14 = 14;
  localparam th_myfunc_55_15 = 15;
  localparam th_myfunc_55_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_55 <= th_myfunc_55_init;
      _th_myfunc_55_called <= 0;
      _th_myfunc_55_tid_600 <= 0;
      _th_myfunc_55_tid_601 <= 0;
      _th_myfunc_55_time_602 <= 0;
      _th_myfunc_55_i_603 <= 0;
      _th_myfunc_55___604 <= 0;
    end else begin
      case(th_myfunc_55)
        th_myfunc_55_init: begin
          if(_th_myfunc_start[55] && (th_blink == 10)) begin
            _th_myfunc_55_called <= 1;
          end 
          if(_th_myfunc_start[55] && (th_blink == 10)) begin
            _th_myfunc_55_tid_600 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[55]) begin
            th_myfunc_55 <= th_myfunc_55_1;
          end 
        end
        th_myfunc_55_1: begin
          _th_myfunc_55_tid_601 <= _th_myfunc_55_tid_600;
          th_myfunc_55 <= th_myfunc_55_2;
        end
        th_myfunc_55_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 55)) begin
            th_myfunc_55 <= th_myfunc_55_3;
          end 
        end
        th_myfunc_55_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 55))) begin
            th_myfunc_55 <= th_myfunc_55_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 55)) begin
            th_myfunc_55 <= th_myfunc_55_4;
          end 
        end
        th_myfunc_55_4: begin
          $display("Thread %d Lock", _th_myfunc_55_tid_601);
          th_myfunc_55 <= th_myfunc_55_5;
        end
        th_myfunc_55_5: begin
          _th_myfunc_55_time_602 <= sw;
          th_myfunc_55 <= th_myfunc_55_6;
        end
        th_myfunc_55_6: begin
          _th_myfunc_55_i_603 <= 0;
          th_myfunc_55 <= th_myfunc_55_7;
        end
        th_myfunc_55_7: begin
          if(_th_myfunc_55_i_603 < _th_myfunc_55_time_602) begin
            th_myfunc_55 <= th_myfunc_55_8;
          end else begin
            th_myfunc_55 <= th_myfunc_55_12;
          end
        end
        th_myfunc_55_8: begin
          _th_myfunc_55___604 <= 0;
          th_myfunc_55 <= th_myfunc_55_9;
        end
        th_myfunc_55_9: begin
          if(_th_myfunc_55___604 < 1024) begin
            th_myfunc_55 <= th_myfunc_55_10;
          end else begin
            th_myfunc_55 <= th_myfunc_55_11;
          end
        end
        th_myfunc_55_10: begin
          _th_myfunc_55___604 <= _th_myfunc_55___604 + 1;
          th_myfunc_55 <= th_myfunc_55_9;
        end
        th_myfunc_55_11: begin
          _th_myfunc_55_i_603 <= _th_myfunc_55_i_603 + 1;
          th_myfunc_55 <= th_myfunc_55_7;
        end
        th_myfunc_55_12: begin
          th_myfunc_55 <= th_myfunc_55_13;
        end
        th_myfunc_55_13: begin
          $display("Thread %d count = %d", _th_myfunc_55_tid_601, count);
          th_myfunc_55 <= th_myfunc_55_14;
        end
        th_myfunc_55_14: begin
          th_myfunc_55 <= th_myfunc_55_15;
        end
        th_myfunc_55_15: begin
          $display("Thread %d Unlock", _th_myfunc_55_tid_601);
          th_myfunc_55 <= th_myfunc_55_16;
        end
        th_myfunc_55_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 55)) begin
            _th_myfunc_55_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 55)) begin
            th_myfunc_55 <= th_myfunc_55_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_56_1 = 1;
  localparam th_myfunc_56_2 = 2;
  localparam th_myfunc_56_3 = 3;
  localparam th_myfunc_56_4 = 4;
  localparam th_myfunc_56_5 = 5;
  localparam th_myfunc_56_6 = 6;
  localparam th_myfunc_56_7 = 7;
  localparam th_myfunc_56_8 = 8;
  localparam th_myfunc_56_9 = 9;
  localparam th_myfunc_56_10 = 10;
  localparam th_myfunc_56_11 = 11;
  localparam th_myfunc_56_12 = 12;
  localparam th_myfunc_56_13 = 13;
  localparam th_myfunc_56_14 = 14;
  localparam th_myfunc_56_15 = 15;
  localparam th_myfunc_56_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_56 <= th_myfunc_56_init;
      _th_myfunc_56_called <= 0;
      _th_myfunc_56_tid_605 <= 0;
      _th_myfunc_56_tid_606 <= 0;
      _th_myfunc_56_time_607 <= 0;
      _th_myfunc_56_i_608 <= 0;
      _th_myfunc_56___609 <= 0;
    end else begin
      case(th_myfunc_56)
        th_myfunc_56_init: begin
          if(_th_myfunc_start[56] && (th_blink == 10)) begin
            _th_myfunc_56_called <= 1;
          end 
          if(_th_myfunc_start[56] && (th_blink == 10)) begin
            _th_myfunc_56_tid_605 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[56]) begin
            th_myfunc_56 <= th_myfunc_56_1;
          end 
        end
        th_myfunc_56_1: begin
          _th_myfunc_56_tid_606 <= _th_myfunc_56_tid_605;
          th_myfunc_56 <= th_myfunc_56_2;
        end
        th_myfunc_56_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 56)) begin
            th_myfunc_56 <= th_myfunc_56_3;
          end 
        end
        th_myfunc_56_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 56))) begin
            th_myfunc_56 <= th_myfunc_56_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 56)) begin
            th_myfunc_56 <= th_myfunc_56_4;
          end 
        end
        th_myfunc_56_4: begin
          $display("Thread %d Lock", _th_myfunc_56_tid_606);
          th_myfunc_56 <= th_myfunc_56_5;
        end
        th_myfunc_56_5: begin
          _th_myfunc_56_time_607 <= sw;
          th_myfunc_56 <= th_myfunc_56_6;
        end
        th_myfunc_56_6: begin
          _th_myfunc_56_i_608 <= 0;
          th_myfunc_56 <= th_myfunc_56_7;
        end
        th_myfunc_56_7: begin
          if(_th_myfunc_56_i_608 < _th_myfunc_56_time_607) begin
            th_myfunc_56 <= th_myfunc_56_8;
          end else begin
            th_myfunc_56 <= th_myfunc_56_12;
          end
        end
        th_myfunc_56_8: begin
          _th_myfunc_56___609 <= 0;
          th_myfunc_56 <= th_myfunc_56_9;
        end
        th_myfunc_56_9: begin
          if(_th_myfunc_56___609 < 1024) begin
            th_myfunc_56 <= th_myfunc_56_10;
          end else begin
            th_myfunc_56 <= th_myfunc_56_11;
          end
        end
        th_myfunc_56_10: begin
          _th_myfunc_56___609 <= _th_myfunc_56___609 + 1;
          th_myfunc_56 <= th_myfunc_56_9;
        end
        th_myfunc_56_11: begin
          _th_myfunc_56_i_608 <= _th_myfunc_56_i_608 + 1;
          th_myfunc_56 <= th_myfunc_56_7;
        end
        th_myfunc_56_12: begin
          th_myfunc_56 <= th_myfunc_56_13;
        end
        th_myfunc_56_13: begin
          $display("Thread %d count = %d", _th_myfunc_56_tid_606, count);
          th_myfunc_56 <= th_myfunc_56_14;
        end
        th_myfunc_56_14: begin
          th_myfunc_56 <= th_myfunc_56_15;
        end
        th_myfunc_56_15: begin
          $display("Thread %d Unlock", _th_myfunc_56_tid_606);
          th_myfunc_56 <= th_myfunc_56_16;
        end
        th_myfunc_56_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 56)) begin
            _th_myfunc_56_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 56)) begin
            th_myfunc_56 <= th_myfunc_56_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_57_1 = 1;
  localparam th_myfunc_57_2 = 2;
  localparam th_myfunc_57_3 = 3;
  localparam th_myfunc_57_4 = 4;
  localparam th_myfunc_57_5 = 5;
  localparam th_myfunc_57_6 = 6;
  localparam th_myfunc_57_7 = 7;
  localparam th_myfunc_57_8 = 8;
  localparam th_myfunc_57_9 = 9;
  localparam th_myfunc_57_10 = 10;
  localparam th_myfunc_57_11 = 11;
  localparam th_myfunc_57_12 = 12;
  localparam th_myfunc_57_13 = 13;
  localparam th_myfunc_57_14 = 14;
  localparam th_myfunc_57_15 = 15;
  localparam th_myfunc_57_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_57 <= th_myfunc_57_init;
      _th_myfunc_57_called <= 0;
      _th_myfunc_57_tid_610 <= 0;
      _th_myfunc_57_tid_611 <= 0;
      _th_myfunc_57_time_612 <= 0;
      _th_myfunc_57_i_613 <= 0;
      _th_myfunc_57___614 <= 0;
    end else begin
      case(th_myfunc_57)
        th_myfunc_57_init: begin
          if(_th_myfunc_start[57] && (th_blink == 10)) begin
            _th_myfunc_57_called <= 1;
          end 
          if(_th_myfunc_start[57] && (th_blink == 10)) begin
            _th_myfunc_57_tid_610 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[57]) begin
            th_myfunc_57 <= th_myfunc_57_1;
          end 
        end
        th_myfunc_57_1: begin
          _th_myfunc_57_tid_611 <= _th_myfunc_57_tid_610;
          th_myfunc_57 <= th_myfunc_57_2;
        end
        th_myfunc_57_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 57)) begin
            th_myfunc_57 <= th_myfunc_57_3;
          end 
        end
        th_myfunc_57_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 57))) begin
            th_myfunc_57 <= th_myfunc_57_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 57)) begin
            th_myfunc_57 <= th_myfunc_57_4;
          end 
        end
        th_myfunc_57_4: begin
          $display("Thread %d Lock", _th_myfunc_57_tid_611);
          th_myfunc_57 <= th_myfunc_57_5;
        end
        th_myfunc_57_5: begin
          _th_myfunc_57_time_612 <= sw;
          th_myfunc_57 <= th_myfunc_57_6;
        end
        th_myfunc_57_6: begin
          _th_myfunc_57_i_613 <= 0;
          th_myfunc_57 <= th_myfunc_57_7;
        end
        th_myfunc_57_7: begin
          if(_th_myfunc_57_i_613 < _th_myfunc_57_time_612) begin
            th_myfunc_57 <= th_myfunc_57_8;
          end else begin
            th_myfunc_57 <= th_myfunc_57_12;
          end
        end
        th_myfunc_57_8: begin
          _th_myfunc_57___614 <= 0;
          th_myfunc_57 <= th_myfunc_57_9;
        end
        th_myfunc_57_9: begin
          if(_th_myfunc_57___614 < 1024) begin
            th_myfunc_57 <= th_myfunc_57_10;
          end else begin
            th_myfunc_57 <= th_myfunc_57_11;
          end
        end
        th_myfunc_57_10: begin
          _th_myfunc_57___614 <= _th_myfunc_57___614 + 1;
          th_myfunc_57 <= th_myfunc_57_9;
        end
        th_myfunc_57_11: begin
          _th_myfunc_57_i_613 <= _th_myfunc_57_i_613 + 1;
          th_myfunc_57 <= th_myfunc_57_7;
        end
        th_myfunc_57_12: begin
          th_myfunc_57 <= th_myfunc_57_13;
        end
        th_myfunc_57_13: begin
          $display("Thread %d count = %d", _th_myfunc_57_tid_611, count);
          th_myfunc_57 <= th_myfunc_57_14;
        end
        th_myfunc_57_14: begin
          th_myfunc_57 <= th_myfunc_57_15;
        end
        th_myfunc_57_15: begin
          $display("Thread %d Unlock", _th_myfunc_57_tid_611);
          th_myfunc_57 <= th_myfunc_57_16;
        end
        th_myfunc_57_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 57)) begin
            _th_myfunc_57_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 57)) begin
            th_myfunc_57 <= th_myfunc_57_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_58_1 = 1;
  localparam th_myfunc_58_2 = 2;
  localparam th_myfunc_58_3 = 3;
  localparam th_myfunc_58_4 = 4;
  localparam th_myfunc_58_5 = 5;
  localparam th_myfunc_58_6 = 6;
  localparam th_myfunc_58_7 = 7;
  localparam th_myfunc_58_8 = 8;
  localparam th_myfunc_58_9 = 9;
  localparam th_myfunc_58_10 = 10;
  localparam th_myfunc_58_11 = 11;
  localparam th_myfunc_58_12 = 12;
  localparam th_myfunc_58_13 = 13;
  localparam th_myfunc_58_14 = 14;
  localparam th_myfunc_58_15 = 15;
  localparam th_myfunc_58_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_58 <= th_myfunc_58_init;
      _th_myfunc_58_called <= 0;
      _th_myfunc_58_tid_615 <= 0;
      _th_myfunc_58_tid_616 <= 0;
      _th_myfunc_58_time_617 <= 0;
      _th_myfunc_58_i_618 <= 0;
      _th_myfunc_58___619 <= 0;
    end else begin
      case(th_myfunc_58)
        th_myfunc_58_init: begin
          if(_th_myfunc_start[58] && (th_blink == 10)) begin
            _th_myfunc_58_called <= 1;
          end 
          if(_th_myfunc_start[58] && (th_blink == 10)) begin
            _th_myfunc_58_tid_615 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[58]) begin
            th_myfunc_58 <= th_myfunc_58_1;
          end 
        end
        th_myfunc_58_1: begin
          _th_myfunc_58_tid_616 <= _th_myfunc_58_tid_615;
          th_myfunc_58 <= th_myfunc_58_2;
        end
        th_myfunc_58_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 58)) begin
            th_myfunc_58 <= th_myfunc_58_3;
          end 
        end
        th_myfunc_58_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 58))) begin
            th_myfunc_58 <= th_myfunc_58_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 58)) begin
            th_myfunc_58 <= th_myfunc_58_4;
          end 
        end
        th_myfunc_58_4: begin
          $display("Thread %d Lock", _th_myfunc_58_tid_616);
          th_myfunc_58 <= th_myfunc_58_5;
        end
        th_myfunc_58_5: begin
          _th_myfunc_58_time_617 <= sw;
          th_myfunc_58 <= th_myfunc_58_6;
        end
        th_myfunc_58_6: begin
          _th_myfunc_58_i_618 <= 0;
          th_myfunc_58 <= th_myfunc_58_7;
        end
        th_myfunc_58_7: begin
          if(_th_myfunc_58_i_618 < _th_myfunc_58_time_617) begin
            th_myfunc_58 <= th_myfunc_58_8;
          end else begin
            th_myfunc_58 <= th_myfunc_58_12;
          end
        end
        th_myfunc_58_8: begin
          _th_myfunc_58___619 <= 0;
          th_myfunc_58 <= th_myfunc_58_9;
        end
        th_myfunc_58_9: begin
          if(_th_myfunc_58___619 < 1024) begin
            th_myfunc_58 <= th_myfunc_58_10;
          end else begin
            th_myfunc_58 <= th_myfunc_58_11;
          end
        end
        th_myfunc_58_10: begin
          _th_myfunc_58___619 <= _th_myfunc_58___619 + 1;
          th_myfunc_58 <= th_myfunc_58_9;
        end
        th_myfunc_58_11: begin
          _th_myfunc_58_i_618 <= _th_myfunc_58_i_618 + 1;
          th_myfunc_58 <= th_myfunc_58_7;
        end
        th_myfunc_58_12: begin
          th_myfunc_58 <= th_myfunc_58_13;
        end
        th_myfunc_58_13: begin
          $display("Thread %d count = %d", _th_myfunc_58_tid_616, count);
          th_myfunc_58 <= th_myfunc_58_14;
        end
        th_myfunc_58_14: begin
          th_myfunc_58 <= th_myfunc_58_15;
        end
        th_myfunc_58_15: begin
          $display("Thread %d Unlock", _th_myfunc_58_tid_616);
          th_myfunc_58 <= th_myfunc_58_16;
        end
        th_myfunc_58_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 58)) begin
            _th_myfunc_58_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 58)) begin
            th_myfunc_58 <= th_myfunc_58_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_59_1 = 1;
  localparam th_myfunc_59_2 = 2;
  localparam th_myfunc_59_3 = 3;
  localparam th_myfunc_59_4 = 4;
  localparam th_myfunc_59_5 = 5;
  localparam th_myfunc_59_6 = 6;
  localparam th_myfunc_59_7 = 7;
  localparam th_myfunc_59_8 = 8;
  localparam th_myfunc_59_9 = 9;
  localparam th_myfunc_59_10 = 10;
  localparam th_myfunc_59_11 = 11;
  localparam th_myfunc_59_12 = 12;
  localparam th_myfunc_59_13 = 13;
  localparam th_myfunc_59_14 = 14;
  localparam th_myfunc_59_15 = 15;
  localparam th_myfunc_59_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_59 <= th_myfunc_59_init;
      _th_myfunc_59_called <= 0;
      _th_myfunc_59_tid_620 <= 0;
      _th_myfunc_59_tid_621 <= 0;
      _th_myfunc_59_time_622 <= 0;
      _th_myfunc_59_i_623 <= 0;
      _th_myfunc_59___624 <= 0;
    end else begin
      case(th_myfunc_59)
        th_myfunc_59_init: begin
          if(_th_myfunc_start[59] && (th_blink == 10)) begin
            _th_myfunc_59_called <= 1;
          end 
          if(_th_myfunc_start[59] && (th_blink == 10)) begin
            _th_myfunc_59_tid_620 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[59]) begin
            th_myfunc_59 <= th_myfunc_59_1;
          end 
        end
        th_myfunc_59_1: begin
          _th_myfunc_59_tid_621 <= _th_myfunc_59_tid_620;
          th_myfunc_59 <= th_myfunc_59_2;
        end
        th_myfunc_59_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 59)) begin
            th_myfunc_59 <= th_myfunc_59_3;
          end 
        end
        th_myfunc_59_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 59))) begin
            th_myfunc_59 <= th_myfunc_59_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 59)) begin
            th_myfunc_59 <= th_myfunc_59_4;
          end 
        end
        th_myfunc_59_4: begin
          $display("Thread %d Lock", _th_myfunc_59_tid_621);
          th_myfunc_59 <= th_myfunc_59_5;
        end
        th_myfunc_59_5: begin
          _th_myfunc_59_time_622 <= sw;
          th_myfunc_59 <= th_myfunc_59_6;
        end
        th_myfunc_59_6: begin
          _th_myfunc_59_i_623 <= 0;
          th_myfunc_59 <= th_myfunc_59_7;
        end
        th_myfunc_59_7: begin
          if(_th_myfunc_59_i_623 < _th_myfunc_59_time_622) begin
            th_myfunc_59 <= th_myfunc_59_8;
          end else begin
            th_myfunc_59 <= th_myfunc_59_12;
          end
        end
        th_myfunc_59_8: begin
          _th_myfunc_59___624 <= 0;
          th_myfunc_59 <= th_myfunc_59_9;
        end
        th_myfunc_59_9: begin
          if(_th_myfunc_59___624 < 1024) begin
            th_myfunc_59 <= th_myfunc_59_10;
          end else begin
            th_myfunc_59 <= th_myfunc_59_11;
          end
        end
        th_myfunc_59_10: begin
          _th_myfunc_59___624 <= _th_myfunc_59___624 + 1;
          th_myfunc_59 <= th_myfunc_59_9;
        end
        th_myfunc_59_11: begin
          _th_myfunc_59_i_623 <= _th_myfunc_59_i_623 + 1;
          th_myfunc_59 <= th_myfunc_59_7;
        end
        th_myfunc_59_12: begin
          th_myfunc_59 <= th_myfunc_59_13;
        end
        th_myfunc_59_13: begin
          $display("Thread %d count = %d", _th_myfunc_59_tid_621, count);
          th_myfunc_59 <= th_myfunc_59_14;
        end
        th_myfunc_59_14: begin
          th_myfunc_59 <= th_myfunc_59_15;
        end
        th_myfunc_59_15: begin
          $display("Thread %d Unlock", _th_myfunc_59_tid_621);
          th_myfunc_59 <= th_myfunc_59_16;
        end
        th_myfunc_59_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 59)) begin
            _th_myfunc_59_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 59)) begin
            th_myfunc_59 <= th_myfunc_59_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_60_1 = 1;
  localparam th_myfunc_60_2 = 2;
  localparam th_myfunc_60_3 = 3;
  localparam th_myfunc_60_4 = 4;
  localparam th_myfunc_60_5 = 5;
  localparam th_myfunc_60_6 = 6;
  localparam th_myfunc_60_7 = 7;
  localparam th_myfunc_60_8 = 8;
  localparam th_myfunc_60_9 = 9;
  localparam th_myfunc_60_10 = 10;
  localparam th_myfunc_60_11 = 11;
  localparam th_myfunc_60_12 = 12;
  localparam th_myfunc_60_13 = 13;
  localparam th_myfunc_60_14 = 14;
  localparam th_myfunc_60_15 = 15;
  localparam th_myfunc_60_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_60 <= th_myfunc_60_init;
      _th_myfunc_60_called <= 0;
      _th_myfunc_60_tid_625 <= 0;
      _th_myfunc_60_tid_626 <= 0;
      _th_myfunc_60_time_627 <= 0;
      _th_myfunc_60_i_628 <= 0;
      _th_myfunc_60___629 <= 0;
    end else begin
      case(th_myfunc_60)
        th_myfunc_60_init: begin
          if(_th_myfunc_start[60] && (th_blink == 10)) begin
            _th_myfunc_60_called <= 1;
          end 
          if(_th_myfunc_start[60] && (th_blink == 10)) begin
            _th_myfunc_60_tid_625 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[60]) begin
            th_myfunc_60 <= th_myfunc_60_1;
          end 
        end
        th_myfunc_60_1: begin
          _th_myfunc_60_tid_626 <= _th_myfunc_60_tid_625;
          th_myfunc_60 <= th_myfunc_60_2;
        end
        th_myfunc_60_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 60)) begin
            th_myfunc_60 <= th_myfunc_60_3;
          end 
        end
        th_myfunc_60_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 60))) begin
            th_myfunc_60 <= th_myfunc_60_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 60)) begin
            th_myfunc_60 <= th_myfunc_60_4;
          end 
        end
        th_myfunc_60_4: begin
          $display("Thread %d Lock", _th_myfunc_60_tid_626);
          th_myfunc_60 <= th_myfunc_60_5;
        end
        th_myfunc_60_5: begin
          _th_myfunc_60_time_627 <= sw;
          th_myfunc_60 <= th_myfunc_60_6;
        end
        th_myfunc_60_6: begin
          _th_myfunc_60_i_628 <= 0;
          th_myfunc_60 <= th_myfunc_60_7;
        end
        th_myfunc_60_7: begin
          if(_th_myfunc_60_i_628 < _th_myfunc_60_time_627) begin
            th_myfunc_60 <= th_myfunc_60_8;
          end else begin
            th_myfunc_60 <= th_myfunc_60_12;
          end
        end
        th_myfunc_60_8: begin
          _th_myfunc_60___629 <= 0;
          th_myfunc_60 <= th_myfunc_60_9;
        end
        th_myfunc_60_9: begin
          if(_th_myfunc_60___629 < 1024) begin
            th_myfunc_60 <= th_myfunc_60_10;
          end else begin
            th_myfunc_60 <= th_myfunc_60_11;
          end
        end
        th_myfunc_60_10: begin
          _th_myfunc_60___629 <= _th_myfunc_60___629 + 1;
          th_myfunc_60 <= th_myfunc_60_9;
        end
        th_myfunc_60_11: begin
          _th_myfunc_60_i_628 <= _th_myfunc_60_i_628 + 1;
          th_myfunc_60 <= th_myfunc_60_7;
        end
        th_myfunc_60_12: begin
          th_myfunc_60 <= th_myfunc_60_13;
        end
        th_myfunc_60_13: begin
          $display("Thread %d count = %d", _th_myfunc_60_tid_626, count);
          th_myfunc_60 <= th_myfunc_60_14;
        end
        th_myfunc_60_14: begin
          th_myfunc_60 <= th_myfunc_60_15;
        end
        th_myfunc_60_15: begin
          $display("Thread %d Unlock", _th_myfunc_60_tid_626);
          th_myfunc_60 <= th_myfunc_60_16;
        end
        th_myfunc_60_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 60)) begin
            _th_myfunc_60_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 60)) begin
            th_myfunc_60 <= th_myfunc_60_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_61_1 = 1;
  localparam th_myfunc_61_2 = 2;
  localparam th_myfunc_61_3 = 3;
  localparam th_myfunc_61_4 = 4;
  localparam th_myfunc_61_5 = 5;
  localparam th_myfunc_61_6 = 6;
  localparam th_myfunc_61_7 = 7;
  localparam th_myfunc_61_8 = 8;
  localparam th_myfunc_61_9 = 9;
  localparam th_myfunc_61_10 = 10;
  localparam th_myfunc_61_11 = 11;
  localparam th_myfunc_61_12 = 12;
  localparam th_myfunc_61_13 = 13;
  localparam th_myfunc_61_14 = 14;
  localparam th_myfunc_61_15 = 15;
  localparam th_myfunc_61_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_61 <= th_myfunc_61_init;
      _th_myfunc_61_called <= 0;
      _th_myfunc_61_tid_630 <= 0;
      _th_myfunc_61_tid_631 <= 0;
      _th_myfunc_61_time_632 <= 0;
      _th_myfunc_61_i_633 <= 0;
      _th_myfunc_61___634 <= 0;
    end else begin
      case(th_myfunc_61)
        th_myfunc_61_init: begin
          if(_th_myfunc_start[61] && (th_blink == 10)) begin
            _th_myfunc_61_called <= 1;
          end 
          if(_th_myfunc_start[61] && (th_blink == 10)) begin
            _th_myfunc_61_tid_630 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[61]) begin
            th_myfunc_61 <= th_myfunc_61_1;
          end 
        end
        th_myfunc_61_1: begin
          _th_myfunc_61_tid_631 <= _th_myfunc_61_tid_630;
          th_myfunc_61 <= th_myfunc_61_2;
        end
        th_myfunc_61_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 61)) begin
            th_myfunc_61 <= th_myfunc_61_3;
          end 
        end
        th_myfunc_61_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 61))) begin
            th_myfunc_61 <= th_myfunc_61_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 61)) begin
            th_myfunc_61 <= th_myfunc_61_4;
          end 
        end
        th_myfunc_61_4: begin
          $display("Thread %d Lock", _th_myfunc_61_tid_631);
          th_myfunc_61 <= th_myfunc_61_5;
        end
        th_myfunc_61_5: begin
          _th_myfunc_61_time_632 <= sw;
          th_myfunc_61 <= th_myfunc_61_6;
        end
        th_myfunc_61_6: begin
          _th_myfunc_61_i_633 <= 0;
          th_myfunc_61 <= th_myfunc_61_7;
        end
        th_myfunc_61_7: begin
          if(_th_myfunc_61_i_633 < _th_myfunc_61_time_632) begin
            th_myfunc_61 <= th_myfunc_61_8;
          end else begin
            th_myfunc_61 <= th_myfunc_61_12;
          end
        end
        th_myfunc_61_8: begin
          _th_myfunc_61___634 <= 0;
          th_myfunc_61 <= th_myfunc_61_9;
        end
        th_myfunc_61_9: begin
          if(_th_myfunc_61___634 < 1024) begin
            th_myfunc_61 <= th_myfunc_61_10;
          end else begin
            th_myfunc_61 <= th_myfunc_61_11;
          end
        end
        th_myfunc_61_10: begin
          _th_myfunc_61___634 <= _th_myfunc_61___634 + 1;
          th_myfunc_61 <= th_myfunc_61_9;
        end
        th_myfunc_61_11: begin
          _th_myfunc_61_i_633 <= _th_myfunc_61_i_633 + 1;
          th_myfunc_61 <= th_myfunc_61_7;
        end
        th_myfunc_61_12: begin
          th_myfunc_61 <= th_myfunc_61_13;
        end
        th_myfunc_61_13: begin
          $display("Thread %d count = %d", _th_myfunc_61_tid_631, count);
          th_myfunc_61 <= th_myfunc_61_14;
        end
        th_myfunc_61_14: begin
          th_myfunc_61 <= th_myfunc_61_15;
        end
        th_myfunc_61_15: begin
          $display("Thread %d Unlock", _th_myfunc_61_tid_631);
          th_myfunc_61 <= th_myfunc_61_16;
        end
        th_myfunc_61_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 61)) begin
            _th_myfunc_61_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 61)) begin
            th_myfunc_61 <= th_myfunc_61_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_62_1 = 1;
  localparam th_myfunc_62_2 = 2;
  localparam th_myfunc_62_3 = 3;
  localparam th_myfunc_62_4 = 4;
  localparam th_myfunc_62_5 = 5;
  localparam th_myfunc_62_6 = 6;
  localparam th_myfunc_62_7 = 7;
  localparam th_myfunc_62_8 = 8;
  localparam th_myfunc_62_9 = 9;
  localparam th_myfunc_62_10 = 10;
  localparam th_myfunc_62_11 = 11;
  localparam th_myfunc_62_12 = 12;
  localparam th_myfunc_62_13 = 13;
  localparam th_myfunc_62_14 = 14;
  localparam th_myfunc_62_15 = 15;
  localparam th_myfunc_62_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_62 <= th_myfunc_62_init;
      _th_myfunc_62_called <= 0;
      _th_myfunc_62_tid_635 <= 0;
      _th_myfunc_62_tid_636 <= 0;
      _th_myfunc_62_time_637 <= 0;
      _th_myfunc_62_i_638 <= 0;
      _th_myfunc_62___639 <= 0;
    end else begin
      case(th_myfunc_62)
        th_myfunc_62_init: begin
          if(_th_myfunc_start[62] && (th_blink == 10)) begin
            _th_myfunc_62_called <= 1;
          end 
          if(_th_myfunc_start[62] && (th_blink == 10)) begin
            _th_myfunc_62_tid_635 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[62]) begin
            th_myfunc_62 <= th_myfunc_62_1;
          end 
        end
        th_myfunc_62_1: begin
          _th_myfunc_62_tid_636 <= _th_myfunc_62_tid_635;
          th_myfunc_62 <= th_myfunc_62_2;
        end
        th_myfunc_62_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 62)) begin
            th_myfunc_62 <= th_myfunc_62_3;
          end 
        end
        th_myfunc_62_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 62))) begin
            th_myfunc_62 <= th_myfunc_62_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 62)) begin
            th_myfunc_62 <= th_myfunc_62_4;
          end 
        end
        th_myfunc_62_4: begin
          $display("Thread %d Lock", _th_myfunc_62_tid_636);
          th_myfunc_62 <= th_myfunc_62_5;
        end
        th_myfunc_62_5: begin
          _th_myfunc_62_time_637 <= sw;
          th_myfunc_62 <= th_myfunc_62_6;
        end
        th_myfunc_62_6: begin
          _th_myfunc_62_i_638 <= 0;
          th_myfunc_62 <= th_myfunc_62_7;
        end
        th_myfunc_62_7: begin
          if(_th_myfunc_62_i_638 < _th_myfunc_62_time_637) begin
            th_myfunc_62 <= th_myfunc_62_8;
          end else begin
            th_myfunc_62 <= th_myfunc_62_12;
          end
        end
        th_myfunc_62_8: begin
          _th_myfunc_62___639 <= 0;
          th_myfunc_62 <= th_myfunc_62_9;
        end
        th_myfunc_62_9: begin
          if(_th_myfunc_62___639 < 1024) begin
            th_myfunc_62 <= th_myfunc_62_10;
          end else begin
            th_myfunc_62 <= th_myfunc_62_11;
          end
        end
        th_myfunc_62_10: begin
          _th_myfunc_62___639 <= _th_myfunc_62___639 + 1;
          th_myfunc_62 <= th_myfunc_62_9;
        end
        th_myfunc_62_11: begin
          _th_myfunc_62_i_638 <= _th_myfunc_62_i_638 + 1;
          th_myfunc_62 <= th_myfunc_62_7;
        end
        th_myfunc_62_12: begin
          th_myfunc_62 <= th_myfunc_62_13;
        end
        th_myfunc_62_13: begin
          $display("Thread %d count = %d", _th_myfunc_62_tid_636, count);
          th_myfunc_62 <= th_myfunc_62_14;
        end
        th_myfunc_62_14: begin
          th_myfunc_62 <= th_myfunc_62_15;
        end
        th_myfunc_62_15: begin
          $display("Thread %d Unlock", _th_myfunc_62_tid_636);
          th_myfunc_62 <= th_myfunc_62_16;
        end
        th_myfunc_62_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 62)) begin
            _th_myfunc_62_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 62)) begin
            th_myfunc_62 <= th_myfunc_62_init;
          end 
        end
      endcase
    end
  end

  localparam th_myfunc_63_1 = 1;
  localparam th_myfunc_63_2 = 2;
  localparam th_myfunc_63_3 = 3;
  localparam th_myfunc_63_4 = 4;
  localparam th_myfunc_63_5 = 5;
  localparam th_myfunc_63_6 = 6;
  localparam th_myfunc_63_7 = 7;
  localparam th_myfunc_63_8 = 8;
  localparam th_myfunc_63_9 = 9;
  localparam th_myfunc_63_10 = 10;
  localparam th_myfunc_63_11 = 11;
  localparam th_myfunc_63_12 = 12;
  localparam th_myfunc_63_13 = 13;
  localparam th_myfunc_63_14 = 14;
  localparam th_myfunc_63_15 = 15;
  localparam th_myfunc_63_16 = 16;

  always @(posedge CLK) begin
    if(RST) begin
      th_myfunc_63 <= th_myfunc_63_init;
      _th_myfunc_63_called <= 0;
      _th_myfunc_63_tid_640 <= 0;
      _th_myfunc_63_tid_641 <= 0;
      _th_myfunc_63_time_642 <= 0;
      _th_myfunc_63_i_643 <= 0;
      _th_myfunc_63___644 <= 0;
    end else begin
      case(th_myfunc_63)
        th_myfunc_63_init: begin
          if(_th_myfunc_start[63] && (th_blink == 10)) begin
            _th_myfunc_63_called <= 1;
          end 
          if(_th_myfunc_start[63] && (th_blink == 10)) begin
            _th_myfunc_63_tid_640 <= _th_blink_tid_324;
          end 
          if((th_blink == 10) && _th_myfunc_start[63]) begin
            th_myfunc_63 <= th_myfunc_63_1;
          end 
        end
        th_myfunc_63_1: begin
          _th_myfunc_63_tid_641 <= _th_myfunc_63_tid_640;
          th_myfunc_63 <= th_myfunc_63_2;
        end
        th_myfunc_63_2: begin
          if(!_mymutex_lock_reg || (_mymutex_lock_id == 63)) begin
            th_myfunc_63 <= th_myfunc_63_3;
          end 
        end
        th_myfunc_63_3: begin
          if(!(_mymutex_lock_reg && (_mymutex_lock_id == 63))) begin
            th_myfunc_63 <= th_myfunc_63_2;
          end 
          if(_mymutex_lock_reg && (_mymutex_lock_id == 63)) begin
            th_myfunc_63 <= th_myfunc_63_4;
          end 
        end
        th_myfunc_63_4: begin
          $display("Thread %d Lock", _th_myfunc_63_tid_641);
          th_myfunc_63 <= th_myfunc_63_5;
        end
        th_myfunc_63_5: begin
          _th_myfunc_63_time_642 <= sw;
          th_myfunc_63 <= th_myfunc_63_6;
        end
        th_myfunc_63_6: begin
          _th_myfunc_63_i_643 <= 0;
          th_myfunc_63 <= th_myfunc_63_7;
        end
        th_myfunc_63_7: begin
          if(_th_myfunc_63_i_643 < _th_myfunc_63_time_642) begin
            th_myfunc_63 <= th_myfunc_63_8;
          end else begin
            th_myfunc_63 <= th_myfunc_63_12;
          end
        end
        th_myfunc_63_8: begin
          _th_myfunc_63___644 <= 0;
          th_myfunc_63 <= th_myfunc_63_9;
        end
        th_myfunc_63_9: begin
          if(_th_myfunc_63___644 < 1024) begin
            th_myfunc_63 <= th_myfunc_63_10;
          end else begin
            th_myfunc_63 <= th_myfunc_63_11;
          end
        end
        th_myfunc_63_10: begin
          _th_myfunc_63___644 <= _th_myfunc_63___644 + 1;
          th_myfunc_63 <= th_myfunc_63_9;
        end
        th_myfunc_63_11: begin
          _th_myfunc_63_i_643 <= _th_myfunc_63_i_643 + 1;
          th_myfunc_63 <= th_myfunc_63_7;
        end
        th_myfunc_63_12: begin
          th_myfunc_63 <= th_myfunc_63_13;
        end
        th_myfunc_63_13: begin
          $display("Thread %d count = %d", _th_myfunc_63_tid_641, count);
          th_myfunc_63 <= th_myfunc_63_14;
        end
        th_myfunc_63_14: begin
          th_myfunc_63 <= th_myfunc_63_15;
        end
        th_myfunc_63_15: begin
          $display("Thread %d Unlock", _th_myfunc_63_tid_641);
          th_myfunc_63 <= th_myfunc_63_16;
        end
        th_myfunc_63_16: begin
          if((th_blink == 19) && (_th_blink_tid_324 == 63)) begin
            _th_myfunc_63_called <= 0;
          end 
          if((th_blink == 19) && (_th_blink_tid_324 == 63)) begin
            th_myfunc_63 <= th_myfunc_63_init;
          end 
        end
      endcase
    end
  end


endmodule

